��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8FΡ��'�N$4b<9^���_.x.�S�}��_�wd�rV9Mz	kb�X]!��:J�#�7�{r��x���:ό���Ȱ�2y/r��m�\�R$�<�V�1Y ��\?;W^|�bAj������h�W<j4�U�e�c�ދ�c�k�1�xix�`J�_f�2�	�ӊ�Y�������-�#����R�9]#�G�QӠ��
�N�< ��/F�+*��?<��i�/����b���X*�ꂖ���c �c����Ҭ�rsoEAC�XZ�M[��������}21�N/'S�2��b� eM�x��44�hVk�
����*6	���ҡ���㛜�
��>�VCޗ��9@�ܴM~�����~���:�[>�!����W	)T�F³�.�sA�Z��R�a����F��S:YB0:�;��Ť��27Xaϙ*);���%r�(!d5cbj�!/Tל'�N�!�w5��f�_ࢇHڊ�U���W�q��)����b"���bM��T��m����7~�.�<!�o�0��`�ˎT�˼�c���&��;��Ў��<���ƞ��s��X�r�Y�����/a>��_�w����9i�#\����h�c0�b�\]Θ�%`�@] �:s���m�d��Z�s����F�f͜��p&GqC����ι�L|�P^L�&!Aw��x�9U\�+�f;�jI�(��� 4W9Lru?�F��'a������N~���B@M��bf�9I"ei�j�ySe��r�o��g��qP��&p��M�����(qK����4;B�y�>׮��f}T�"�|��f�
G��՗$��`p��Z.��T�F\4��hD���x��O������ū��D�'�N(cQR@M����饷���a&��3����~�~V]�"N����{O.���ת<}�pgU��Y[bЍϠ�g�_�̿��&�WA��܄�Rv���c� ���0t֛ӄ@��2ʅ1�AR�t�@�g�,dP�w-�"����5� ŷ�u ��ш�AF�|�:(�T�{�P/	��a����VJ몢n❬�_d�3� F��x��0�b3� r�q�]"If�Q�L��A��l�rX��1�򕑘�����G󍹭�!�V1���B��?ھ����)DG��󀼶��D-�Ɠx��;�y���z~�F����0S��>v��᷼-�xiq���I�Q͊DK^�'���xW�(�h�����E�<�6z+w}�`uz�ީ���tP��vO�(��C�!�������v���w��{��[�]���,}�(Fr��;z�ȐT+
)M9�'���@���|���-A�â%�`����<� -�.�b������N��|�8t=/1������m4(jP�`�{��L�Z[�Q��D�9���!�сJ��h��6������In���t��F��D襴X�,q2Y6x�T��T9���|b���K�k�j�P��A��2�%I�������<f�d�N3l�V���QѠ�a�V�����m]����T�S0���Cү0^�J!V|!M�T����f�L��p��g͟�TA�Hx�l�B�k�ԋrf �;�#6� �6��f3-3� }ҚZ��E����Y�U3`@0� ���7e�7�d�G꛷�v�ل�6�a�����{
��!-g�l�@WG�-Љ �ؾa�{��LU �����(��K�`�S�ݵ���O�O^��tDF�:@�	�����،N�38.b8ے[��P)�Ͳ��3����ЕRe��ԍ[ϱiP%��:*�=$Q����B4�k�PI�.ŵ�O*[��j���)��!x��m>94�a��� �UE-�������A�'�~Py�ྵ��Pj�ߟ��]'���5�������r�m,t;�����^�3d_��n�b���G�ZDa�<4�
�Ee:��b�奜�7�=��1�l��+��`�+\�Ê=�<ǐ�F�9I7a����	�k0П���Z8��AmY�.+��%$g�P�?�������H��a��M�� ����c-����9�$	��u2 0�n��7EXsk�h?��eْ<|�Ѹw���#�+p����C9�5�á�{��q}�}��st����݂6R��¨Gd#�ѷ$Ws���Zѫ�bب�Ч�N�YԞ�mw��E!7���.��3�b���*��~@�6JN8�>K� \&�o��Y<"Є1!�-V�cae�����w��UR{�'���#�c�:?+U����������3@��o[���q���D�Y�#�ZBPJ�^������__g�f	���}�>�I�Q��Y:�?V����2��s{����*�s�i"��Fnp�3��_��gi���6K���)� �zN\����-���Yo�x�����.���4��dE`��L���lH�"n�E��Kxm�K׶C{� (��Zw�Yg=|LIU[sc>�X)�,q�P��#�A�$�!�~T4<Z�,iS*����M���q"���4@w#�!|�f�����af]���f�%Ϋt\��A�|���̄��R����į���%7��&�����M��L!�x�K
���x+�-�𑫻�&����(���� ��5������I��(\1���25���H��`Anw��e����Yig��ky.i�
��7&��'x���n�]G�c��E��A5k0��P�'���l�m)V3�Sz3hlV�g�����ұ#��O �v����N���-##�V3D/;�8�H�չ�e�}��a�I*��Ƶ6`��EȋZzE�D+;|E�p1�jX���ɗ��t�$��u��Ω��x�<�k���	�����X�b��&��tI�Oވ���\�Z����� ױ��Q?�Jp$���xp�E ���}3��e�۠�}}���(�Q�O�	Y�������?�+ln���Py���_��O.�%�n��uBE+(�x����Oa��݇�.7q�J��Ȍ�k���20�r����/�A���q	��v�ŏ����rE�l�*ߑ�!��C����aJ�b.�܀y#M�*���}Q�nނwy����=��R�wp� I�`�řz�fz&Cل��A^3q���#���c�`��|�7�;**�|�&=e�/<�D��l)�.>�kJ���B8R*�!
�j�g��$�yTD��r�ҩ��)��m���B��X�򦕱'�9~�5��_7��B%�G�م��d��j;5���73�^�����7�g��!�:��hP�4��߉��#Os�Z�lC�m��Z H4���DS�Ă���Ƥ5�G�����&̶O'S�׉f�L]B�{������#�wg0g���e�"  �my���Du� ;�҈�xI�o�%�A�\A!ڣ����).��v����ۘ�R�TBV>��Ws?���|�5Ӽ9k4�]�0�F,H'S!�fem=^J��0W��C�i����zl+�D;�p�q����m�E����X���A�b�	Lq�݄ġ���Z9,ȋ��%>���a�
-��x�ۉ�-��a P�X�w�l$2��ӫ�Qo{j>�x�-�s%boe%�Y���E�آgG�ƨ�����=�ݰ 5����ԅ����d�p9;֩)6���H���=���X�/pA���0�,��"u?Y�z�6�d�}Bfe��'X�l5�F5�k����f�z�k@��F拴��A2���L�B������u� �sT���L��v?Y� ܜPA���pN��g8j����=`��{9G�������,�1�@()ѡv�"�rG��'|���J�aQs I[���843�8FCU�nD3���� ,R�&7�k�븬��/�v�#�~uXd���%��-8I9D��7B�SF��`�_�ϋ�;Vq�CIg��;�0˲7:C�r`�7=U�#;�JI@�wq���kL��S�կ��ZK��&�#�����Ek[F���u�% �}��t�w#U���<�~�ՈN�N;���������o���gva2��8�(�ؾ�]�E,����lҼ�{�*��� ��;%*� 0����D�����#���xs����r3����Z$C�A�-�Q~�,$�#Ki���L��I��(��(<�����L]���l�|�&��_�-��e	�Ae`�?Nl^�a;�PodKp_��&E�1ً��kP�Eʰ���$��d��ϣz�0��5mY�h ~�u���k�Wy�
�K����kuxM��{�=�A������'�UHCKȌ@�^-^!n��PWϨ��.�	��� 0�)&+2"L�V굍��z��-�x�����o�Dӎ�0���+�%ߘc�k!�j�B�6�������L�֭�&�k� �9̺ZR�����eIQ�"]��H#�;ٻ�`4�/�����[&�t���=����6 ����<�Q
�>��@d�Δ�YjZ��Ů���?'�?_o0��CH�*%dfٲ�ۂI�Pb�����j�j��sc���kG�V��th2�Md�S�#�w��O�9���	�Bcg+���iWHAI���K�9Cz�&og�������R��O�dA���p�[�uv�Mӳ��y�t� ˝�E���������"L�72F<�	e9��5!&����u�I� V�CXc��:��o,Bj�!���H��qģ�5��M_r�8�#d��>oЩ!*dW�"J_� o�p��5�C�a2�ݾS�w5k_��sp�A�ߵ
�#�߾�+�}}wu�33�5BF���8�忰{s3���4Jr�`�t�'�*a#�mĤ��F��a���[< ��0fU]7U�vL��y��?���G�N�x�T�Sk��[[��E�ͬ{�~_����>�����W^(,�:g�	~�;��R�
��Ҥxj�)�!���YWi~[&����FpɊ�e_�4e���cR��c$��Q��]�+<��HuCv�>
���mR�L�"o	b�))�X����$$�>ɤ��������r�,��q�UG�[C�Q����C��75רtޚ��:�����qD��:�3�dO�$hm�!��G�/�����0z8)$���ȉ!5 .+DQ P4F!z�A��k-T=\P�J/�Ϣ��3˩�B�k�DA�r�+��~�~m�!#Ozp���e��I`���_���7�ї4�"�4��=7#,��,�� ��9g�h�"v;ˆ_dǯ �db�Ͻ��b��ŸI�:s$ �de�I���������}�xdV*N|����� H�#�+�(t;�+
li-�{Z��u�l�v�G��þ��|yE�S9�p���|��~p���?'6�F��Fjn>2�~vI�b=���;2�^��,h��c=~��(�~�O�K�7���*P��F�ǖ7���D��P|ZV���:��&foQp�#�-T��i4&8y�U�� ;�Y �=Y�����f"�|/��e���� L�>����^�$-Hּ��9琬=��z�k��.�T�����p33�d�ᝪ�Sb�Xh���(xAv�8���d�v�Zp.���w)�w��۶�G?ymW�Lz򖅒�i��{����2:��lG�2�AL�z#�d��*e2�1�Px��q��)$��31������Ɗt)��~ρ�JS �z'"(���)[�¾��MS�?	��0�?�����3�����9��ǒ-"³�y�4�R|�w�Nw$yyX@*��P[��#������ LG�j�_$�g���-A�M��3$�����pO%?�ǯβ����;9�r_�%�}���N�މc���n�i�ߝXi����'�y��Fb���k�'��L�cP����R�{�[B�*~\�:�`�ۙ�c�Z��P�:l%{��9�����ka����^�x?[o�' ��ĮG6��W��I[o���&�
�"vd5|�^���Ey�ay�$��Q��y��[*�HR�PW��۵QN��W�/qp1� $Y�&�����U[+E�� �����=0�k��#�k٘j`�������C�Ęlű������O����������Z��d$?�Ҕ$F-�ޡ�?���%G��$�z�V)�+�0�tƘ�'�����ܰpy�O젽O���Q�~�<%���=؞����SL�}�p�ݜ���.����ăpP�#EW$6 ��s	Ȑ�D�$�´V,�M����	��z��Fj���Rǂ�!�O#z�ݥ��ٯ�|���'gx��7�.)J�==4�k$hp�PhL�@=!��4ɛ�E�a�4��B�{w{޿�E�J��N(#�$l�T����p�R� h��"��f�y�9�m�����o��������2E��y�������_^
�H$,H�kP��3�5����U.;oI�Y��E�ș�Vח~����y:ʎ��M��G�o�G�"�{���� -��95�j��(�������$�����(L���t<��ɍ
�2�F�]g3:@ـQI�� c���bo|��K2jT��,��+�ow c�%�~PL0�7�8ƝC��:��Ռ�.�/7�ƃc��u�c�eg��y��! Ϙ�#��_n(ï��;h����z������z?i}�1}�;�q �M��$�!�Ov/�� p{�/!z�����J�g�=��ׂk$=������硼�ob:I� $�׏�ϸYԭ���p��pњ�$���mr=��XH� ����zV fδ�H玔�m>M�ؿi����ž��� ,�-���-qHY�L�<�ߩ�9V�8�i�����+�}���2$���j�/�ӝ�Z��I<i�P-�~b��J��If��ȕ�	`�vXMD:*��x�� P�{��1�1,/��	�g�������>�ċ�I��~���)԰[�7�3:���;j�{��჌�n�r��.�[�m|pz� ���яcIF8dv5����E�{	8�p�{_B��{Z�P��^�}�ѨN���x��ļ;/A��<~2~>vG|@q�s��z��X@��ɐ�pN�;�_��<��ݛ��76.$�QF����[��=��"vnzP���,�w++��T���t�T�$�~MK�6a��������]��̇#�ɝ�U/Y��yGW�����]Y�3&au�<���L.�)�4A:����|5�AI�� �Kkrz6����#6`��>aZaj�����0
����]Q*.�����6��}�S�>����bo�u�,Y�ɹ��ʍ��ĿG|k�v��f��Vs��1�t�#9�K���|� ��6�մ��tR�D���P'd)�R석�7)<������?#���Q�?i=�|��p'����$����$�����w{���k�\Һ6|#�H�tҮ[ꚕ�es��ʓ��CP�g� ���	��$�1QJ�^�f[;�B �	�y:��}���1�G�e����Fj.�d��Id3L]4�q�Z����f�d�w4e�	bFH��߮� �R���J�Hף(d��ɶ��͑a�8�o��ۓ-

�kx��Ly�'��'3�hU�D<VXj>3�W��L���'�W9�V�Y�q��x3��A��3�,wc�Dӳ�������s.���Vz-a�>�������]��7�����(��v���7��g �\�T'�O),{�ZC*���h��v�o�G|b	�G�
���!��$#�SD�T���K������/����'`�n��Wf��o{�c�$NɗK�i(�v(����z�V:��l*%��q�\�d�-wpCy���:7\#�B���q�S6�G�f�Fu�>���1���rY�*�lPN$P�<S@�� Dy㧏7�KNL��_-O��qI�c�.�u��B}�B'HP��t|w�4���7�A�\���Q^���> ["��S��Q���"���`�h�J�+p�y6��_UĢ.9{h��#ؗަL��&� � ��ˀ�XR�h�H��������V�z��yۧ�<����o\O`'�*>�ϐ��PX�}>���G���g��#��:�)t$p�2�ٍ�����H��6��A<� ��E�Ȋ֞�n֟'3&���o��9U�e�Df\�� ��#U���u<A�+�aI���|�	��L�����P��0~���.R�6.\�|߳��8��C�|����y�/��7��lC`���:�>�X:��\�&����Y�eR�45l�V�?{�O����߁ʐ 
ל��.�:�����
��G*q�>Jo����c/rgw�A��ٙF6u��K%P!�n������Y1�d1>kw%�}�BbÒ� fS��������D��w��v���hi|���o�܍(s��L=.���P���r���]�^��2�>���zI���݌��;R�Y��JK�0��mS�:F"��%��0�!Q3�����u�	�j`W�KZ�:W�\ۙ	n"�R4[�v���b���qM���[_�S�tL�ꅎʂ�����o���͔���`hi�;��ΒGA.���y]`kMd�n)��r�YM��]�$��-S�(\_Jw;�XW��Å^E ϥnc�kp?g$�k�ro\�}��.V��֞_��Rf��J{@���KF}ㅸ`�0�����G��M�R&a!%��n�g�:�����?Ȁ�^7Ál��:�� ��s�yN�Ŵ!{"	�/  �`�
؛���c�:&�����9�g�i'ۤ�)d��s��T���$��ǬC$ݜ�Y$쨉�H%�Ӫ�n��p����!_ݫ�u��Fs8��@�YF9��H16�>�$�e��O��@���-x�;`�XfD{�"�ݶ�[s��EI�;}d9`�)��R~�o�+��ҫ٣_?[-ߤa(i���; '�\�sQ_z �lA�I+ᰟ���9w�6쌟+�Y��k�u��	�u���D$ʧĠ��}��\j�fj�BI����R����^`����W!��sk�($ANT���+ܗ

w��)ɡ����fɁ��9��6��c��ј��9��\g9��z�艒. �\P����̽Hs���}7WC��qL���U�#O���HA���J���#��3C��%��\(e��d���FfK��Y�I��@#�6�(��o��o�M���~m�e����oo�����f���f>����V3������+��ހNt#:�(Ü5[�3� *n����0=�:�\aH���`�����[H��ϛ�ߎVd6ƭUP��J�+��3��Bcn��cZ/�4yۻ���1���� �������`�:Y��2,ӛ��*A�s}u`����s� 2N��!���O�5�G�_�x���b%ut��/�A'՛��	)�0=���� G��F��?�!.�.S35��M?M+��b���Y��$�Cd��f��pNG�TpF�z�3�ܷ��q�PHx!|+�#X�UA�H�R�m�m��g�k8�Ak��(W��T#+ �Ő6Y��Ɗ��<;�Rt":&���Ќ�|RHe����'&P1ZK3^�g q�p�6a��,ǟ�rmx<���S*4����D�7�!�W`�%}1t�o1M�o��56���sK��4Yԥ�Z��;l��_�.�&��;`$C�����t�������`K\ͬ�E�=��7 ���ÅO���"fs1Y��w��j2N���g#�IG�����T�oj�}R�O%զ�p�Ql~!�,�����S�Ӥ4�IQR������l�A��Zpe�P���O��O�}��L��,	�C������3]V�B�V�D���$6��$��ef��q��.ڭ`*��V��X}r�㔘�$�9k�Rr��:�����5^c�ЍdZ�+v��Z	9��J��R����)�=�ot�~�t6G+4Ra
�i��C.����`����)��U�
^�X�ؿ~�����_[��Q(�� �R��0� �1�t��'y�A��P����I�GЦP@7O��^�#��L�q���^Vr���^�1'��9�୤�7�����x/��F`[|y��Y�T�>TG��c�'5u{�3ca���Yr�e��i����bvADzuwt���[s+��� �3�$��g�b c�2��;��q�
N�vq�$gH��v`ٙn�{g~�
�f��z�\�,��h>'ʠ��3qBN)����1W�U\q&X�p-��X�h�%��ǐƎB�������]��'��TA:�m�/�=��20B} �FO�s�W�2�l�w��A|����ȟ�:�����M@.�Qx���mn�e~lN	܉�կ'"<�ᠥ.5 �,!u\R�������FN�PoG�x�npAЍ��RHc���=ܬ�5%�ݎ�=:�~����C���)@$�6N4[��� H��9�2<߸	�����Ջ�`7b��L��و���#�y�#���:�cv�^���+�?��_�O���N�x�5���,���s��8u�Hs���^�}�\�q��
�C3��tJ{��V? �or��2�
Ӝ'��Go�xPR��Ĺ��Ś:3��*�� �.]�D�k�,�*qK=�I��8�D�֊�;�K���"PW�%����>��P::�g@*a��o�@�B
�:K/4�sq��ͬ��|)OQ�Xv��.h�[�[�����n.Y��w�D�u�����׿={V0{�i|MD��,��SH��n>��:���n��bw-����L\�K�/mpZ��c��؊{
}ԙ)�Tg�Hg���$<;�V���:?\I ��J�8�h�ʽ% L�O=�-��ڳ �o��`��.e#�p�����k�x��S�|���6����߄�����3�?Q�3Vg�b�qMc�Y��<�8"��C�-�#){��i�H`�������a�H"w.�+Qh��֜-��8��q��r�v�`�i@ d�O�/��z�ih�ߟ��@�-3"�(P�s���#2�����g�0F�m�"����
�*�m��(���8���R�~��χM���C�N��3���d�W5ل�v�fw�;����6�k��Oib�{ۿ�8�<���L�-QB��x�W�pi{�	w�й$�v��rH�ћ�]�����.]T/�3�H]�M����C
*[Υ�H3���K��t]mz�v��7�S�°"��])pp�񘩤&�Xm`J��j[.�����~�ό���r���zL>ew��'�P�6\�pi�j^N�x�K�Z9�h�	c�H�sG��$O���m`�v���9�AV|�ƳUC�zp=i��p��w���k�z�P0p��P.L�Љ�Q�+mRޱb�Θ�,y᩼�Β^!t8	,k���y.�d�2P�P�I��q��m�#�7�U"��![_V7�͈10JT�u���#ߎ��L�-&�&�6��7��j�!��_*b-w�����{F��실�V�c�Q�k|�0 �NC����W �!�^}9u��Q�qP@��I!�Ԟ>���n��v%���
�#].b_��g�؂��z�G�n��;�Jdߌ`0� ���4�讞��
��$#��U�&��zk�fVWY"`	x��A-�	�����@���;���	�ԣ�Dȣ��m7�x�m�X�9��;�:��t�ٵm���om}��6�mNW����[+f�Iӊ̙i��U��c�Z}ՏU&l�zɬ�bu�l�MǛ��>��4��-M᪥��]sb�J��c	Ť����%3U�d��t ��k�H $�hH���!t����Q\WR��lo���h��d�e��;�O��#���e�$��9�>�dU��O�?~��kF�w+��)�8�%�G����?;��_>�w�F�<>>��6�=�X9��ׇ���oG��ٚ�v{w6�uGr��آ��?8	��5
�9��t6�\�(����69$3���zoh�w�e|�
�C��d�HN�ላ��6�t�,vt�1���| ����KM�Κ4@Тe��}5���Y�e7p�bO��]�t��k�s9����\�z��ʏ"�*@(�mT>�	�`�<@��h�@)O�ice�C"F�Jp{��0�͹��-�	JΟ�(^j-еP�v_��S �7�_��8#^��`a�}�Ƞv��Q��OhF��YͶ�Pרt�s������\2�c��Z5�k�h�U ��k�3��>��U��LH/J�U�\�P�TT�A@��T�?yy��
��ݎ��*\K%�ƈ�+>X�Sˮ�pK����gt�#^o�O��U�����n���E@ P�Bz��L����Z�?��	r.|E���h}�ؠZtQf�j�p�Ϯ[�@�бב�������M�"o�
���c��m-��� d�4\P�n����p�(�$.�~�Ob�&���@_(�+.L�t(I\ۊLf�W"=>¼��G���&y���ݬL�Uf���e�Bd��� t/��KAs�ߚ�&� �v�c�1:��aF$췜2��{0 �Cpq�2&cT��-r$*�
,t���֭���<�]������熞<Fm�S0��2���rbFo4��R�F��`�F��vh��QK��w�&�;�Ĳ�G�M�-����=6���pKYc��4��#�C���Ҭ�ؑ]X���=�'�g�V���1{KsW9b�݀l+2T���M�<颌�hy�Nk�`kT��6��}靚�'���X�FP�z���J����OĹ�,�Y&�މ�
��e��?//�� �4> �(Q��[❪gPzH�ﳀ@ͅ���.��t,7��J o����*N:�E�d�s�6��	i0�b|0(tsՉ�T8����`2�� �Q���+$Z����C��!���u�Mq��0����)a‴ɬ�|��g�4�Y�R���bn��x��#�s�a��	
����Z�;ʑp1���7�C�^�){qi�Zl�6j��$uL��:�NI��Iرy۞�`B��)�0Ը6���I��	��Yߢ@eUx��ݯ��jRI�^յ�:3l鐅�����j�z(5�N�Lf�r���GO��Bxi*�\�p�A��1\>� Y;qJ�2�%��a�⑝����0"�OFP��Qj��8]�4�R8�m�B�����a
�O�`"P����B5i�)|��l�Gˆj��N�+)�8��Ƅ ���fP�

��ta$�(�Zd�E�'�U+_��&'��%K9�ӗ�z\��vU��&\V�*���4���D���G��px\*N��=�m����b����/���n�v1�k+��Io�����#�r�A~8,o^	�#U�Sq����ss��4����J�II�$$�r���(w]�@1���ɭ�����~1\-�sۅ�Ƌ`-��w�d����$*C�Cq�uU�m����f<'^�p�.�-D_!d���ĳ�+�k/v��'�q��my��+���>H�ef�XAp��7;|�N������:�Ȱ��x���H�<�G"�����uG3o��č7ܭ�Xݭ\7U����%�7�|	�#�`h�B�쉍��Bi�x�/&G4���G98Z�J2�㷲H���I��I��^�*0�2@s�`&�MrR6�V՘N:9B;_۠�|m�O$�·����ǳ�ǴPL=5��?��4_��c	��~^�e�+5s��]p���=f]��X�v�a�\=أ��fN3m|�r8�'|F��O)�%
]���G�et6�t�=�!ᜧLN� x<�-�����C}FU*�9
���~��y|�[,b����?w	2��v��_��*�Y�l���6�X*ٓ��Hm��o�H��<R�6�P���.F��%�J��j��)�6h���PQ��n([|�EjZ�7��Gt�l�����go�^��O(Au�޿<�N��>	E؅@?�J��8�����Q���)8�fy�b�gi%�a��Y>W=�Y@5n�)�"3N�����^^vP�!��[�Po���	s��eS�p]�Zm�~{�js�VġK���b�
s9n�����F)���\��nl����4�{�EO=z����	<d�:uU�=o��=�����S�n�N���N��iܘ�٭0e,8Y�1k�7���m�~��j� ���+�@Q�V�+1�ǯ�6k����}�PSD���3�D���IE:d�p�Z���\���41��60�7��~�$��=9��M�O�{��3rG��[�Z�:ش�� >e�l�=>nAt:z?�u,��*�S�z��}�zwn�1X�r�M�������S/������Z���~c���R�l����	7��YeP��MG�~{�)'S3�IZ�bU���T������]��D}����֠Q�Xy��o��^�ZL�����!߳=lr5EWP��s"pZr�H&v�AP�sC!I\�߈��*ߘ\�i� 43d��t"W�� C;��מ=��!w�Q�&l��q�9�~��#�h�$L�ɠ�L�E�a���a<�v��ǭ�y��͝��x}$�X~O��󝤃��S:<�c~^)�gM���,� ����x�'kU����p�*;w>pvY�i���ݲ(p0>��Ww���η7�	2�.��!�3�miwUIg�Go�4!��)>���G�q����h��j?��'N@�@�ۉ!��n�=K٢�eA[���?�c8��O���1f���Vz�8
�L�t�o&�/*�L�m�Kw�S\�q��?���8^��1�IƾD��R�9X}X�d/�W8�K�}���,���wH&ϧ�
�!h��.�{-�fYc�������w��&�Vj^}�ҥ|�$���Yy�۪�x�
0���Pwx�(��~�Z\FS�o���x�@���X6J�m޳L�A��I~Q��c�3�T���_9:���~�*�;x���yP+N�7�ۮ��|5��l�	�dZ�I��K)��� �F( B�;t�W[r_~HMQ<�~/�<�O�$Z�\MȬ��6U�M�"��$����o�ے�Eo����`�/V{b[��E%(�ѱ�N�iT/ǒ�2��թ0�o�BdT?��z��$f�,��Z����!5����9#��a[��F�.FU�hy��hwƶ��Qu�#evNڧ;���fb��T��9!n�`5��]�� nƄg�Gd�5^$gO?=I�Z�S!T���/�b6&�8�ڪ��@�]�j�?QD��{o��
1&�!Uv�6}la�;��t��� Y�=�#��G\��sl�A�8�n��}��>̑�� 	��B'{�&E����q�;�#)�	��� ���B%y�ڵ\�]|�\Hح��r8|8�r@ nN��%3�?�����'&xAu�Fd��;r,D/LR6���3 l�z_a5F��4����PW[���s��߄j�e�a�6?�����S[��u5�"{ �u�J�Z_ѕ�I:��F)�����%���-,oUt�%����B����ډ�o`��4�v�\�W������I�n�A����:�����"��BG�H�*�D�`��wS�Q�"�r����zD:X�d�ѹ:Z�M�,QE>B���j#p������Z
o�J��.$�Ŋ�*�X:f����6!�/�-R�����Ua/���� ��l�ʇ�LU$1��l2�[�_��j�|J�;���z��6�EE��k]�.�G�F6�h�Ƒ0�ɳ�L�H+b���<^db#�(%>�yт�X�����) ��W���\�2��+5�C�B��Կ��`��mҷ�7;f1,g�{:�*=8Ʒ\y#i'�o)���CU;�f���cL2��)���ŠL@1tsЙ.���w!�����^Juh��`��������^07�Y��s*鶇:����ɉvx"��l��[�n�Ү�ˡ6���YG��n l_��癝����#���`w�E_��("E���&�0p�\u7e�s(�E��B��xu�>�`#��	��?FdOuяr���Ċ��e��X��ӌ̚lK�%���P���朌m�.܋�I�:��p[^`�ի+�cޕ�,0b���g~�mZ4kM0ܸ�(��K����hյ�mT]~�ꢪ� U�Znn�g���7]��}�����dps?ȪY%�h�d!:t࿵Q�#X:R��вx��.N8�b^�������+�"�3l��o�d������k�|>Ѷ}h+:���[p��s��Z*�`�:�����i�N3L=�D�+��.p�E�����IV7���Z�Q^~�*�N�Q�� ���_(��K��yf�Z��/PB(Ķ����X�u�
f���9�|ϱ	'��)I(�����*���L0����h=�Ӳy�h����t�c>�QA�MYja���d�^��:m���yi�'E���y/�6�];򞯁sq`N�*�}�_%ѯ+�2H�p~�/"f9��))U'�tE������;��M�Ԇ;1�*�0������'üK(*�9����|�t\�Q\@�� ~,�e�Ԧ��F[m��*c���A[�K��y\I_{9��/	����~`�?��\o�t�iۺ>��G�z?��$$j�!B?_�P�sx3�#�T���8Z�怖V
�	\,��xq�	 ,qN",�V�-|��K����[7$eh�nڼ]�D@wnBKք��kҹȟ�M��U��>Ӻ�,��
Z`ه����dz�5���N .(y����I#���ŰҬ���ʈ�ToA�(i����ƭ�σ�/`z�� �*�|�_S-~�s}M�C��(B�	������ٔ�5��n(��(�*n:xM�UY�{5���
T�&kʸ��^��f��ŤV���T�zU��m�P4�cs⎲�n2T�R��K{P:�5�6�FV|��R�˜0�3LM���L_,E5����	�sm"l�����9�`(�.�.j���%a,k;m[��Rh���#,l���55������q*~F���zytdݱ��_����L`�dyFSs�dIԹF��^�7��N���LU�9M�?�F�<�ӽܡ`���VP�[_�N��խ 2Z����DѨ (X��+��蕖k�j�(�:����=ds��pt��yx��	sI�[��9�X�tEg�Y;ij����).]��nܔ����r*�*��$hPvе:�.�Q�����-A�.:�u<�&��ϹjL��j5��"�90F�,��[z_C��<�B/��?��I|�a��9Ǽ|���!8��s�,�Q�� �O�!�8�T�c}�m�8�#W�
��p���.)�΁����C���TK^ k!QֱRX�ʊYx1��S3��A�k�0R����O���Ɠ��"5��q�jP�	�~�[��pV?uXl�s��y�[\��尋�D���2��KED[�t^QӜv?[{y���&�4�nwX�mc�-�M��W����y.���S,��Q0"-W��o��ص[����WsД�.�V�'��s��CtP��E"����DK#j#k�pC i�Ǣ6���9��`RsU��"����=0�=g�vF�X�a� f ���$�;ja��4�1=��(�m����`��7��G	��<�r��czrЀO��]�d�֐l�7���^��r�čޝK��S�;�?<�nD���q���Sn��M�.%#E�f��Z�-F�U�I�qB5��oÌN����J��[�wvyܗP�8HCa憱�F��� ����|��p�u_�dW6��_0c�f�erU���qx���k���#�1J oS!+�O�U�;���aǍ���Nf��?ݮ���OF�xşpװ\��ou�k�^MA7�A��p�����6��1��������Ղ�^�SQnOQ{�s)|�_z"f�M	���|�׃p ͖K�M*�m��ww�g�x�1��M�hH�pR/]g"1H���#�p�����U���\6l��{�x���]J���;А޸Y.�w���-�a�j�*�<��%�{O04�������� 
��� ��I�4�
Ӽ��,ģ�6����h���ޖ¿����������ש�G��O�܎BwN������Vb��3���~�VHBHY�^���KD�휝�9.�J�O}�zG=�QZ����wr�Fe�xܼp?o�п�3��
Y�A�������Y�)��������{V�7�#����2�y�a���_iU�;�4Kz!��8��Ǉ�
�4����P�G��V�	n�x�]�צ-��{�_��ϫ~}i���	O�C������Z��
?��T�%���@H�w3�Z�����7'.�(�A��h|�W�kd}7ӄ�qQ���1c�5���d�AUg��a���+�^K�.�]01	;!��.H��cՠο��.ËWSg���I{�ǈ���f@d*��	 ��\ctk(=��2�A��%G��N��c"��5T�<���}������xr&E�%b���#�A�W�ë���a�=L^�Ƥ���՝��LO�^p5�/��e�:} ڮ��{��ҬNB��3������G�啄����x_7ќ��'{t��"�#�p��0x��	OzG���z�c;e8�ݤ��/�W�?��9���{��|�e���̢�O��i��@U;ۇyNd��]W �\�Pɮ������W���T����VнMn�cѝ`�_�!O5�x P��>E����M"�pVm��5��xB�rzJ`���-�E蜒�f.��n p�Y:l��\��`M���4φ����B�Hq��V,�̓�6����,eGg��!eoظͲ�\������\���Rи����Ղq$�Y����F֘���"QRg&���� H��+�C�HGrhǡPH������ I����YY''ά(X��bR+���L�,΢pl��gա�fs�w�I�#{�1{��	�YP���C�B���4H%����NZ�gc?�MpI�i]�㦏��p�\���;���,��>�5ϵ�m�4�
�F=���$ޣ�����Ҩ����uH��������Q�]�|��`4��׳�=X{�8��ֿ3Ni�6�
��޵���*����;��]�ޠ#�M�/-��ɔ�?��1�S��UṮ}�N�!�v��f��-�` ;.﯈��U�+��产��1�T!��D�<� :9��c��&U����\זA�w����������u!�@���Mj�=*r?qb���(e�#mï��[�^t�nv��J�pV�ҕvT2�|�]�i/:�e[�����h�qٝ�|��Eg��ɝ0.���Ve���_,q���k�+}������v1x������T�ooB�I!�����ְ^�<�w�ԩ��qdn��^��W��TO��!���P
e�Jv8��B�k��	��&��.���̶s�V�Ģ���^"�
-I�����)d$u���r9�������G���.GE'_�m�}�W�vy�h�� 7b��;��L|�4��6����|���j�#�C�'�n_�/�2��9�zF�	B ��~����zܢ�8���qF"�wC�ر��g@F�%�C[��>ɠfn�oeW�,N9W0�+	' �-��90����J��j1>?�LA�������Ew���7Xh#ԍC� ��[�m�Hd��_�?Y�x��ޛ)���	O�^�C��`��#	N��L%+o��NOIRë����\�{�
��@���,I-J�2Oy�K�4A�ʛr����1!p��w��D�X�x ��
�V��L%�s�$QD���â��\��2L�>j�����1�"�4��_,��.[룇D�{ּ�֏t�����n!��Z+{��y�R��T<~�5�>TC�����K]Ǩ�L��Qn2�m4>t��9��;��3۹eQ��4��T}Y��{�7�\�(��U�Lp3"f-���iֱ�؝�3���{��^�.��>ʵ��;��o�� y0�Se���y�:���}#𧻛S��)�?5`T]�>�v�zW|��<�0	��&Y�jY{����!ӷ�7H.־���8�a�-�Vb0�(T{�t{e�����`��Ō�F��#n!E��u}���(�t�!c���6��sl�Z;z��۩���8���?�8W)�2�ĭ�4&�,��#�#>Y�]	f���ѹo|!r<,����r����B*N/�,-�t�,^�]$Y��08���3�%���h�O݇ݭ$aM �!���Sm�Q�kf���ߔ�b����9�0�=x��1�o�Ɩ�#�j{���q�C�E��AG�r�]c6f�L<`UhLC|)��<oO�};l��8aږ�O��n�F��7���|�����[K\ʮ4�9h5k��ܿ7Q�U�� ���YשX�ǒL��]�o����w�u}*�v��4�)��ǟmiGٟ5m�d}䌲(�:lZ֩�m~l؏/�-4�
��DUu��������~�f�"K���e�vkmHY��a�)��kd�W����) �;�#��x�Gd����\�I�x'k�3Q���`\X	�O���WlC+	�A�y{�>[�#�����qtY��kG�ൾl��$���I�T,�V����dڽؖa��E)��(�����EzsJ�U�r�óIءU'����#�o��̼ܐ��o�0
�1z���2L3��7�5z��=�w��ÇI).�Ίj�ꮧsS��A�\�\�����Dw����W�uQ{2N/���S����n�Bև��ŦA��AS�9� M)���ps��zBoИ�r�\�gm�fr��T���Y��*�o$<k�+J�('2�V	�r�w��Nbt���ݔcD�E+�4���B��<��J���G_O63V��:d='C�5�;�`�k-��[�4��.�i(��9Q��j�Of�ddQsk<���3��2�a�s�]ݒ֫0X%J8"4ȒQ��#�L/V\�^WfUU`��@q)LZ�����z��� bu��'n��8������>�����2\GtY��"~]��T�b{���{�(s�����2N `E��K�B���$.�(Z�=������W�������ͤ|>�[����ғ�x�r. 5n�{�:��H*�#I�5ew��'q|j����Dg>�����z1�ܨ$]�v�g0������<�(5w�f�JF��ӣ#����������b�s�� �R',a���U��;����,��f9�����$?�������r�x�cq�����;:���œ�q��$ A͏��~Ĉ���U� 'u+۰T����
���B����m�RN�
�+�� �i��`(�C`�l~�f��^/=�>i��7!|B�����\b��y֞G�cA!|�<�����m}_�y�?˾��ۺ<'�ZM�����*�~��ҏnarJ�|W���C;���q>}�,��p���>SJ��$M��2L���-�P���7��,i���W�#��ƌa��'������6��6=<���D�Z�[kLA��!�ڛT���5�[_!����e����ʀ�0��*"LFʸq�)�e�7y���e�Vk:��9ˎ������D@�/Lr��5
Ѱe��ۺ-�͙U�4��D��5}|��gCI��4ĒF����;�H� �/�������`�c��~[<��vZ��o�*�Vf'v��P�;S�P��>��/����L��Q�b�B�YMy�?08���* �U���)�$F��#;٩:�W��3�����Lp�uzkz:G�ThV���� �΃Q]l�n_�������"�7��V��h�͝+G��Rox/�!�/1)���3a!n̲g�T�6�C~��_7����+���V���e{6(��1�!�lr_[�Q��4��<�3�57��v�X/��� �FW2A�[Q�n�@z��>:w<�&���tc�o�.^:�,�4®R��VߣxZ��0��Y&�i������kS�v�!��Z��ߒj�1>�o��)��ƺ��?Lԩ?��s1�h.��h-�A�=ft+�r�$88�S2b��ZUn���.���s�~�:�"�76¼!�^��L��?�;6!7z��Jd���{yB��	&���YL��c�c�e��^&�@O��Fdv�Ym��?A�C�����+<Ģs�v��.��Y�X"�b�ƊG3���%j!�9Jf�m�n�NF�y��v}�Z���r�nw�ϗ��pn�g�\�����|QU��͂��3lz���ǎ�7Q3�"Z�]l:?�^��q� tV��8	$o�}�6\�Mh1��U�J`��󟶨��w�W����F�]3E� ʹ���GQ�Ū���	6�+���"E�ᕌF}�ل\ �8 � ƣq 'fǙO�6u��m���YTR�w�7�V����x������\�����T�a�l�CC�8�{"'G��!?1�x��DA��y���UL�t�D��Nҝ��*��h2
���@����1���؟g*�$�0�Z� �'��{�H$;�eÇ`��s�/���9�9yx���B<�ٞ<���A��b[��8|�"����i�cC���97��ِ��}\kPZE���$�I'AB�{o'z	����$�Ogό=I��qO�ٯ��1��*��V(�2�֮:<���Ηh]x��E!�������Rl�:����U֠���b��l%2m�x��y�T�`�4��!��˨�ğ^�|Ww����8�!-r�,�G�tV��R���
Z�� �$�M�������֭ �9�L;�6G���;������!Vw�V��	 �����ol&8)��xr�Y�L9NVy����+���F�Tx[�r+r���6�	��Wi&��a�K1��Z�)�ӼҞ�Kr!8�F�E���rW�ʧ�~&e)�M.J��h�p��*Q_7,!o#�J*�������XN��/Ƕ.�cy'�Y;$�?�EdE}7U���Gp
�&���w꾑3nwSR�'���=���|�����TV��Z���>�袠0{,xO���v��?�k:}(���abh�rR�ٌ�.�b�X]՗����(���]�9���&���jҊ��k�Td��q6wՓ��i�/s�K�|w�۞��ŧ�����a�Է��p�a;{E�[tE�  $�L�v ���1}=��J2G�-��X4�y�)���5�'EڔqؙemESύ��� ��αA�t6x�i�v`�?�P�Z姷p	f0����ZU |�x�l6]%c���U��ۛ������'�YP
�^�٥�IU엽�*j� ��Z�;O1J�"aj��d�D4��04�q0���l,e�lݠˢ�G7}u1eq�.O>3�8�V?�} �I��xvx�η�,�ԕ>7���Ȃ&�x��tP�9m��$%V�jyc�)D�c �Z�-��k���_J�Ir����&W��x��� ڮ���O�w�p���d���&�1c�݄�-�AHL2{{�u�y�0���K�0�R�~�L�)�Db/u����zFa�s�u�Ko�現�<�Ъ=��x�a�v?�gp��"��H�����}B2��a�+s7��B����g{���{���Ð�ԋ��QXs�雊��Ma����8�AF�Z�Q��!��T��P������
��Y�DH�*Rk�'��U	ן>�6I&0����ͦ��`���!c�>�J)�����ye�e��ϋ=j�u�s&����"�.��.���#��Z>��β|ߝg��+R�'�8��DV��v�����
^V�j,A���Z6�Z�|�J#�7������D>U6����8�A�0}|S�8�h�6�1T<c��)�qfTV�`5# #h��	د~������s1�$7)vl&���a0�;����@9���H�F:�fW��l�@���}��6��<:��a�5q��枪b[g���0��ֹ�
�o%���� v��r�փ���C�d�U����!�5�n��ÝS0Aໂ�[;A�8
֊��5q���S�u�+�1�،\���L������<��Y}n�V��A��f��|g� �����$� �R>-����j�=Tb��O��A�;�k7#��ł��͊�,����(�kDӡ����`���E�
�d^ ,�|3*a��g%#Gk�м��xōo�=�B2D�]�l! ���y��1�b�]�/�䑪4�}�G]�.�3^�y�B�����Ŭ��UBM����Į�˯��	�����t�4�H�m��{L3�K~�V�憛�z"�c<�����g�ƿ���9vOw*V���Vl7����O6�����D3��+��|�xov�����|�!]���������i����q1�{��)W��8�ʇz莳���@�4��~����\0O;Ԁ)�д�����=�����
��̂�%hp��I�L��Ȟքo�}O4����lM��Ԣ�A���P��#�j���7�{��kI��w<������b��kP��^�\��X��$(.����e6� <��2�i���V��?U�����GH]���v�����ʱ�U@�2fs��HvE�֙UO;���5�Vi8����򥾰�0m���8+T2FST%�f��>e˥ΐ�o4fo�*��3�	߯�Z7 ݥ<�@3}��+����Ƀ���io-�k?�n#`܀S��a���f��ꃸ=�$��a�{,g�?5�#!꯹aj%-Dm%��Mwzu�"����B:�P99�Hm��s���rg�]+؋Bˊ
�y��O]��:�u�5�*�Q&�oݔ]��(�?j�Zn���_Hȶ��P��p�b)6+*`�>f�����0Oe���W˴0�\��8�n%^���r��RpW��yr��O����{!Ud����Fβ���]D���[�p���f�0���y=+�[�撫vɿ۶�L�R#"O�{�ʻ��	�r�����H)��
�?�Qnˡ8�:���&C\;k�?�1�VA�!	��8�hP�F��R����)�I�q�zHd���^K������%80'���Ҳ���S��{/[��k1[*�F�B�ٔ�+�K)�,cr��XG1P�锔�]�IQ}Af�Zk�8�X�:aH���s���ݷ�%���rE��S��L(���uԪӀ0?����� ��7B���⦖C�V��������WQ���K!t52?�"����d���rL�@��\Ի6�윜�M9��~������A{���A�\k�d{�e�J)Ľb�`�""	��V�< ĆE����235HI(�����E%>:�_�|t�2�+B�h�A<�����?�^P�W����wi��O��4u�h%
�E)MQ�����)�c��5M�G�t4n����#�P�)D��W[s�@F�)Z�ǝ+�����v�i5�R�Ը�n{İ�1��$Qd��6�ow��#[i�oЍ��*�:wj�~9��O�@%�����go�ed�>�k�ʯ��S��Ob����Bq�tHM��4o!��D�U	ڄ5/�9��Z�o��I"sRt��gcx�v1}�W�JM��D$���c%��ϫt�`x�fƮ���1ݷ�$Q�1D���d:��<��QT)K{?�o��IU܁�A4ت��,
�ͅ��Č�	A2�jAeCy\��n�VC��:q����nG��d���	f����{��q�̻<v]Al�PB��$�2��Ʊ��5+��墇��f��C��Q1��}o�^7�ѵY	��p͡�(�(3�c��a)�o_��)_��V��~k���P��N/>%y)�}d&���0��>w�.���;��C�\X
��f����c�;3�J��̳��'�$�wA�`?���p�@�w]E�P�n���tvi-�:3ߜ��O;P�֪��,���8u���H*��-�%�*���n�1��r?.�S	��*Ӷ�5�a!�X�=��E	��8��AaXG�8��������u��i���o�����hu?߀f"Lʮ���˄�����2��`� �N�(Q����˴�G]/t��'
�q[˿�����8J��w�-Vi�R()�fC��!��6����]��/�@�^'�(@T�W�<~j[X�����4�k�^D
�O)��	�XY{���O�T���+�Ŧ|�27�B4-����L���`�3��0A"FX��6�qg�_���%�BJ�U'�[�$�*��Z�ʶ�~I��Df�_�_��o��E�������x�M#r���4s�I~y���HC���ҏ�m��8�ǃ����ĩ��v��� ̱F���9��]G�(��#U��o���H�RA؂�ĝ/����&sEf	�>����8^��M�5�N�`έ�����.�T�:A-c4kÕ�� �&�g����Aselp����g
�[�?�|<�b��y]���;�_J����ȭ�(~�#t;fI��52�8��:���>���,T���9��c��ͬr>P�� �e��R�vB����� ����/%]��<L��R�Q�B�}'\��'F��l�1ݶ�y�N9�����i���A7��w��"�|(�ܝ%wA��C����v��?�+_y�e���.�k�i��v`�gDC�2�П�ܼ��m�x'�W!*p�׺ϴ	��!�rR�p��}��X�Fd��H��eʦ�s?�N�P8}9d����p��o.B�I�2����㰗�@|W�INs\���>>�ܛ�{p3H����LhP��YX��
��z����17��ϴV�'�c7uG�s|� ��i����O�S\�,�'�6�ݚ�R�<(��U�x��G��#����Si��Ѝ��h�)��G��piE��I�^�ϻ����mB	,|Y�8ʀ��lK�A�;�4r��)�uU���N(wYf���&��(�c�{�+F�%џ��v/6�xrw˲�PB��>�=).L;������@N���f�H�UYH��#�1�	�ŉ.O�Lv<k>\`裺�=�N��V�.���S�}�N�[FS�`p�b�ϣ�[�*�S��v-�p�Ɉ�K$13u∌|<�pi��#���q0C���V���P&�͓��4�|�*c�=�bq�Y�b���?5U&B�j�7d�~�pa��n����	����+
-�b��)E;-d�75��P�6����;��_f�ٶ٭�k#�\*�1Zѯ9�l�.v���9ePus�Xx2j D�~����I"83%�8>x��]�x!����j�fk�|8ᚹ�=���!���%e�&.Nx��˓�k�$�d��5u��am ác�`�=B @����6�0|�
^���tӥ��ҿ�{����Ca�;��P2f~� ��ޫ0��II3��� �P j=�rȼ�Ƽ#�꽻�$n�U~���Ԉ��Ӊ���#��ŕX��I��x�?�'�+R�f���DUQ��:��U*�]����B�<�a�cChE�]�pcˣs}��0���	�m.��F2�]R�N9�L�����)a�b@%�pH�W���m��KB+v�n��H^��O;<��Zb�5]<'I������YF!*�ک��m/�C��Bۗ��'�&�1�] ���{8޲j��l��k(ԗŲ�\��U��e�R��cy��%Y�Ȯ��"C��p��Cpn!��?Ve�	폧�f ��A"�`d�>���Nޢ�ƙ�q �Z��H��n����. ��=�5�0�_�d��}���]##���J�㳫B�SW]��������U>M�p3�L(c'hB��vF�y��c��<O��;A����$5��h��VW=���FLF��%�����ĬFڂZj�B�N?�s�7�6�L<։���Q���n�k�R#�I֩n8?���4����J�Q�����[ڙ�鞅9	��#!�u:\7y�
�%�M��q!h�hV�C��9��s)�5+g�R<?�w�i\,@ZB�0F��D��Ɲ5Τ@����y�q�T�u�����Q!�q�� wr��kJ��&&_CZr������A��8E<�W�<f�|�ެ�/��VI��A�-�&�����_�g�(�e���t���U��� ^���}������ 9�(��lDe��dX[�V��#���s��@ʭT�X���G
&�GC�*���t*���5�V�=줉��D�ZQ(���WFD��m���0���"���w��-K>I��LN�3���>�
E�N�l[E\��z��;���N�kB(�-#��������N7����:H���t�����������'ru���ŝ��u�O��z_ �#���w���{J�Z����9��a-;��"���޶�ΠH�cn�w�0�R�T6�1+Xg��ƃ0_K
�D<C�-A|�E��8h��x��]�9(_�}�G)�K�?E���Y�=�>�<��v�П�s�ُՑzM�C��M'�-�t��]�T�0w�A!���k'�4f�<���u^T���lS6���j+���	��_Gt�"&�1d��TW�1��^pk��ŀ�����m�����h����r�?4���S�jYG�&�󨼵�z����ň0�w5E�����o�a�u��ø/�0)$%B�G{zk�?^�z�g:)�A�$M3��`H|sD|\��F�K(��;+nKT�R�\��{^lYc;Ie5��_�jwN�T"^��>YexrK���*M�}M�&��x?��X���,B�H˞�?��!�b�:	r�e�J�@���DO{*֟��y����O���L�*�S�B�{�ҽ��6dw����X�����8!��ĠZ��Y����Bc(�h?�ho�j����g�.D��@� [w>�����_ �_0A���]�T��	G� 6�񶴎��=����Sƅ��b�f��7��7�����[z��܏2+�7�§�Ab?@#� +�^��i?�D<	{��2����/�S�����gH�#Py��C��!��&�淎�6����:#��3Gw�A<�ޥ��
�0��?���7�(KL=<*��M�k�$,l5AK��7GO�{b��oĭ���@�*g�$�a!i�-���A�z#��)��1,ە޵�I�H$4��q�{�����P�WPw�-X���rS
�:�"�y�D룮�3#~]��������z�G���۷J��~6ޛ�!X�0��5���)���Cu���a>D����c��,p��� N�$�)�����(@0�]j#X*�ENG�T��7BQ�-�#_I�ө�h0�&��u/��EFO��H1Y����v	��!A�r_s����Yi��g���;n�4(L�W@9�"�%��\T��rجCJ���6�I�[䠛�o���{�kX2��*qW�f_�0���:�ӛ��4jB����]�0>�o��Z¬����`� �2h�p���͞߁2W����&�6o�g��7��X/$�Ǘ�����2[xN���W��4�P��.5P8A�� ��ٺϠ�V�f������UH��#ʹ=vi qX��&���|ZX�*?�E�&.A�|�0y��:@@��ҭvr�?R�ߡ���Y�����M'{�<����I�YɏN3��8�%=�԰>Oғ�'��)�
ɋF�=�0����ho��DIL2���t�g|�$��|�xn&��$����v�w�^������-?��k�.V��=�H��=�[�(�*U�Z��L�!:�^n/�3Z�LN�P_3y�$h��G������V�;ԡ�25$��NW�a([3�?�ݨL�G��q�[3E�$p��0`Z�(U�Oʤ2n��yJT��$�l��&A������pA�k:�dP���|��	t˸��=6G*����I���*���Ϋ���
':lφ�1�DjckX�˙��PNh<���|Ee�>?�ϑq�+�������cv
����}>{e$B9��~�ҁ�D��[k�Dr\K.�aq��]"�tP���K]��ڌ����@Kϲ��Ŕa�}l�l��/Tq���e�uִ��|~4��]<Q��4y_ߺ�$���2�*��w�
G��c-���;��0���k�9��;�����	��.รي��m{z�ۗjU��8~L��;vv�:.9ې�Ȍ��J�����]��-���\ �YՔ҃+�Ӧ�����A��#_*��;�7(��e��Epp�$j�˒GQ5����l��&N�Xy����=�]+�P�p&�9��Gg��*�a���J_IB�"&6X��x���p�&�?�q�r6�{�ّ3N|�6^bȯ���e���{Ѻ�z��?�-!��1<�Vez�,�ԣ35 m�Z�QP��}��v��/�A�]���5`х	Bn���ٚe����\#m���uH�>h܇�S?��*��#��w�D�ـH�H�i��uf�:���'�Ӆ���$��(2S@-}}�B�p���qx�pX�bHӵ��!8��6Ra��ҒMK���drpH���:	pD��	;qYW��C���^t�a��t`;���)r�r���`|%��{�ҵ��~W�:J6�R��i����7��۳Z@aR\j{Bl�2�`�}�wp�%�)4,��݄�H0sL�
�{�U�eƔ��ҕ(��T�N�Xm&f"������"��;�k�9 �2�D����D������҇��2@4A�1��>%�L(?As�_�>�B=�Q��2G�H���$ Z�����I���O��8_��OlZ�Y�YJ����������|��7��A��Y��?h��[���&������k�KY	5	�1�?��1�C0�Z�A�g���g=;�JW�H��Lc)):�8�9"ε���4A�e#��Sg��0�2vU�V������?��f�]�t�y�9H��O�����|��=��J1�I�wO��Z���:�u�doB��L������/'Z=ҭ��/%�$[�5���^
�F�K�R� �4���ň�ѯ���q���y��F���F�w�Ne]&�> �B�7�P�*��O���@|�����rd>��:�(h�6�|zd������/!-U�_ȿ�N�$U���:�-[s��I	Le69�of�C9O��:X�+�a��~��K���})�N�M� �	��`��¤�?��q��Xj%��J�#8��z~�w���-�9+�6o�{ �i�AM�u�����>Y�W�^���<ץL�*^,p��#��L�3��1�ۗ��'�ΏPd^9�O��2RP�䉔�	[�/�3
'�,���~Ƌ��|�ս�@C�Ʌ�Tѻ��$��1O9�#�����k��ν�ޯ���uy4����f�#�ZS�tȼ�������DB�L��:���rU|oy��-n�X��$�B�i�*b'�w��E��3�{p��#� �����)��O���0��"r��{��E�vc���8�K�� ���~E�6>Oi�E��~uJ�j��ݹHx[�	�+�`�R?�{\��$xHp��ƒ�0�gü=���HW<��t�4����b�?�؍��!W���Fc�,D$�c�z*���$;f��,�&��(̚��(A��x��F��$nM����	�Wx3���~�A��ǉ0��9S���I��.��+πO8h�B�/��m���LZ�ੵi&OB˨K���;C	}�V��S��h�;�c��j��Ԗ�����F���I�\��WJ�]
��c��9��a�49Q��T��ʠ�ƒ���4���ձr-4c������b ����$4��2.�����u��~��E3��7K�U���S��zhQ)��,�:Q�X�jG��w����˰��	���r�j#L*���{�=,�/�4v��/���	��٘��ʽ�qz~�o�ȠY��-�b�����2_��^lՄ�$E�*�l�TSG��⏵�U�P\����p�[��2��3��j�x=V��A@�0��FnKK���G���0-�_I��>���Z�$\�_�i7e�m�I�AZ�o��4Gћdo�;��#�h��a�,��|4�hU΅��6Y,�R�_�faG�8��F�#��8�����6޹�.~�e�g�������`@γL�G�{�Ji�~^�5��J�%tј  �C<�����:we�c$Z]�P27��A�p�Z��!�>�S����}#�������]��b!�D�κn
�̓.34`������8�G��[� u�r������T9�Y�"!8��3�U����)���C�������T��Nx�4z��{e*��ȼ�6��p��_m��W��	t��8UɬV��/�?Ir�F@�F��)�0�����a���Nǯ����0\ݳ��� zE��e��.�b|[��B� ��f�>(��.N��`�,n�"e(|�{�g�&�9��������5���l片��6f�ݦ˿��H֦���{���C,�Nq����dO�cJ����I�F��HS���һh�]��1A��u+x�dMv��T�>�S͇�����JN�8�|fl=�?���~�8�Og��)�W����p2��w��|%*�F��C���扦_a)��_�k� .���`Ru�q��>/h �S@x>�� �1��S} l =�R�Qj��L�q�q΢+}���0)]m�n����[�1�ߒ�ˤ��ì�qW�_vg�@����a�o���4��yOT"�R����3`4e�c�Pfx��"��PV��%1=�\ ��<VIs�|?��P�AK��8ŷ��b-_3z�Kkc�N�:~�8��p�Q���{״��/���b*��h�դ���T��/�NQn@>@w&^y�c��K�dP�d���y�L-�R�l�n���f�5����chw
$������²�)��j��<���U)@veD��"�.�M���=��A���d�),�C��g0yq�m�|��\��z�n)�:!�Z��<�1\u����
'�oD����@�ɮo�2:*�X�WV!t$||��^?a�Z���}�W�� �®nm�/u��҈,�'R$�DN61��#`�?�4�����|qB.!��Qc38Cj��<UclQ��x��E D�����Ԟ&C�H$=�_P��6?���)k9sFr�$��#������\B�I!�q㵽�{栲ʛ��3��`���ԫ��Ŝ^�7���&���E�̢�˻$)�Vy�g4Ѿ:��6%�S��."G[����G�r��� �Щ�����	��:��0Z8��'�θ^���9����j��1Y���ôq,X�,�>}9�ޙ1`�.���\�>E���<���x�i�-��x������y�9��X�4g�����D�����T	\*�~0�~I�-01�a��-wY�`Fr�A��H%�����U7U�����	��h��E��̴�n�VFL�p�o6U��M�7��־8g��F��g����7�x���;����?S���U����z�p6Y_��u���\Gc�}e$�ީ�y Rd��r�<u��TG.4�W�� �|:�X���T�kK#E��)v����n�|C��J
ZO:��p��I�WS`���  �Go�v��n?�(xe����f\g�@��bW��Q�2��U�'~N�;F������n${=�S^E��x�+�I�	{�cV��e{��7?"� ��MO7W�?��NU��T �")h��>f~�TF�l�97Z��w��wÜ�-�Yv�|Qy�h�2lX���������=B
/꥾Vuv�L�W���|�&<r��
|b/�:R����'* �;''X[ȷ�q�d

ږԝ5��O�1�|+�f[�k��A	��d�y]�vv�"sDNI)9+��OQ/�m�&R�n�&���m�����;�f��b[ \��z�_��\�����k�oR	T,�[f.h� �u�Go�n�et��rA�~�ϹvT5$6���)�4�=(�qw�y���E��Ӕ��2��--e�;����IZ>�( �dS��84r~|�G�=��0*�8�G\=�b>V��Q�⿼h�,*�ՀO���P%�>ֵ������Y�Ն�W�8)G4<m�|L'�2��A��y�0��`��r�ro��<�qʰ�ƚ*6��L7�V�6�ʡ�,E�=!�+��
��rGٿ	@���wSQ���HUC��������:��4j���,��=�&�]��nu�ŭ���% �aPv���)��Ǽ�k�$2yY
�����A�,�HP��8�h�[��Np@�e�����Y���MZ��f�Vv32��M�E�4���]Z��$:���[��=H���j�l����Ϩ"�PD�j���ahT_���s8(��Ag+�_��ķ���m|�~�02Sc�-ۆ��
�i�D�����&\7����0^=�Nmt���XH�@�0�v*:�a�:H��M�6.��쭽�ߊ���x����f����W�y]Y�X
s������@o÷7�j �ww,�1_�9�s��ｴ
Uqo��a���e�V��c2' u��IN�?E����\ZG�N��aц6*/����1AJM�]ט�4o���$��`����W�y�M�k�ի�@�`﷭�L�
�.�E_OG��g����ݠ��l�`y���8v��V�5]�8N���'��i�}d%fY��{�� -E�%Ms��%:����_�Wf �]��n%hb��\A��8t��li�%�C�hn�p�d�%��^>�#�|�D�e�)��a)GK�AjC��`��P���ni�ڦ�CK9ï��9�Ж�:��t�,q]��zl'��5�����{1��Β���׊s�եƚ���Y��VM*��=�>��Oo�R�.���:z�'=�3tF�$,[�<4L�+с~X��%��\�:W��Zd��]\�.���9�&л!	�ھ'��3�]$N�́CJ�3u�I�/�;9���� ����V4��v���"�$s!����֥g��M�Qy�{Ubj&��Cy��c
n��9�%��~<�����?7D�
8C|T9��	�:� ���&�S#L,�f����&H��!"��aĽ�d%����\/E��ޥ��y&�0s��jw@DY�":Yg���*�9dŐm���"I�@ܾ�~�q�����Z@;��_!�F��"�f���/��� P��\���w�*���ǫ�1lc��Q,6�3G�c�&�g+��g�<�������e�G�h�H�ނ� ���P��Pet\j��ffT�/6k��Y	ʢ��4�=+�?tI�t��1z'.z��ٗ$���׸�9iQqL�9���2��At�Ov�mД��
��U℣${[�spP(�?�+��5`�f��"��C��Ƌ8�'^N?!�Ա���4�I��г���P���\q�O���ѧ=�:C7+�4�Hg������_D� ��`��Uzp�����r��n�	�UK�RM4���Wh�"�x��s�6+hrC�	��-r��~�#mI?H��pDI�����ʾ���C
߶��]��j�\6�(���������14r�	�'F��W���̥�y��b [��{��2<K�T�꧇}�۝Q V���Ά �)�9�'�a��f�L^w�j�V��*�H�i���P��5 �FU� vF�m��*#͏�np������@�����U7=|GH4F8Z�t@�Sԇ� V���U[��%������u��>�_t�׻m+����C'	]z�@���r�j�C�Ee�խ l�{U�[%i�c�i���-� g;�8�����>*sFl�^��5�.K¤�cϋ����rn��#�e)�Q�~�}x�+����B�f1��-���H��JT��ȸ��苄<y22S�9���!~CD1�y�b�肆�e���x����.C����3�c��F.��я~�61��<E��%I��R�Љ_�1kެ�hӆj�0�����%��-��c�Ydr}t�,�_�w�V3��{%o���0$���AU ݇T��5蜡'9(.m W~ͷ�ۂ裡*9v_�7ۅ @	�Gx��S��D���L3!��
��G�KwG�c9�i���C�Ѧ&�G�����|�
�&3S��.�z
���9���:�7�I�&�Ui���cCMY^���n��ؤ2�{Ջ�5���0�o���X�+.�g�@�5�D@�_��#�H¾�i�W�;�'���r���ΌkBF ���(t��q���U�{E3U��Εj�jY��ϥ�V���g����3�یPE��w�F*�s�[*d����@�H*W�e���3�t�b�q��?��`Э?�T����E�<>�Ĳ\FM���������\��D���"� Խ��K]�Ի;��fm�;Q����t&�����ۨ��y�z��A�����@C�,�uW����^�l�j�Aɚ�IՀ���u$u�P0���z���CΠ��۬\,�F���^?i0|y�l�}?�ot���2̬I��9y�VCO������� �4S0˘%\���ˤ���q��y��W�Q�ex9�/�`�ji�k=���p�I�p0y!͓�<mՖ��������krS���ج	j�./)[X� ��E�aY=IV!�?&�!���ŧ��ysx�'�6�:o|��6�m�~OK֕l�����i��9~E\T&���y�ӧ�=����!��&S����Ig4X�����k�i�9x5����t���!`?pna6�ɉ�E�.�6���.��o�.S��Y�IK��6��o-�DIa�3o��S<�\@�.����f���9�68�y���u/#-��ԡ�Z�ŵ�`�D��3�P3=GSm��҉� �9��N�w���p�^2յq��^�D���S6|�s	y�`�{���X*�ۡ0�k
����y+C�>��
���i�,Ps��8�j��}�dlU1}�q��3v����&.q����}iBz��jR:X���,e�,�p�xs�;������e~L�7;�|����י�Z6D&1eLD����2��'y�-A��)G���*k�|q$߮�t/Ē�"�ݏr�^��¬��J��&��2�JOgb>����/�ЭbY����q�D��{&E�-:͝[�2K��A�A���z�-99��푔�v�`g�?t�JH���	H�B���(����n�T�aa�lHFV�Dj�������{8$�}Y�;���㣹�jZ�?��'rS�Y����G˕���=��D��������&��cQυ7�d<�:x��K�ki���l��t�8FJ�b�n��6�?�U �*'�O፜K���fޔ&�-dӬ��W���2�HNf��&4��면�K����z[��5�<��jD���ZB�����=�\����QW�W��r6�YX�3��'x��:����X���2R��F�Y�A��F�go�؆:	>9��M�Ԅw )���^a�ӄ*0i�ll����T��U���+��l��kLvZV��Å�l�=�-�P�A��3im��EJ�[NN �"�V�e'��w��۲�܇����79���_j,����:�m��DCt]j
%64�8��\p�-7�3���c���o�ˎ\g����	�(�,�U(L]N��b�X��+�rMir���+�6�Luȇݗ�cz�o�l)���G+��sոn�P�Η`XK|�[~h0��f�A��(�ߝ�#RD��Jw�t��DPP�J�Yo��\;��?����!���"/�����W�����#���T�У4F'��I���3�f�w��+p�hp�� F3�~
Wz3Ҳ�T%���G�ۿLvV��#ںbUAo��n�r�&-�x�gp#mG�|H��A��8����Wэ�=�0����U�]�?�;DT)�8�H�j��y�]�q�������o|����)M��P0X���P�[Lq��8
hG��:�^RC�� ��,���t�޸��}6�<r�A\�̠�^	�%�� ��;�bZ�Ӄ$�%�h(� ֘���l;����|����K\��_.�e�҂��!�h���;z@���9���G�M����^�T��x��1�!{���o����#f��Ma�JOu{+�}�N%�p�h`%���\�k��UsZ���,@�?g"�[��c�^���1p|v���0a���G������_�I��,�]I��/���+�*M���J��$��!dyQ�����lkl�e�Fx�K�X�"�¥��%򺺎����c����j:!�g�r��*u"�"L�Y>R֖�H��/&#�Ge_�Sʹ�"A�96Hv��7�nPn��k���
L�E5��,3��P�p �E؜��I̀aM���v�r{4�'[�J�
�:��-H��������5�����u���V#{��<�����WiU�g��w�O��=� +6H� ��^�ɘn�\�yQ*l,؅�
v#t��C��	kFm�R�*�A�JT!	�۾b�kpڎ`wL
+j��UX�F�Km:���'��sޗ�i���̾9��"h,��� 4lːD5L��ѳ;�n��B�_Aq��Ru.��&v�t�)�W�<a���1q�C��h~����^�Ό_}z� ;�H3�?s�|��`�(iɞ�87��d�����T�6�7��]����5��.xͶ��,.��_�8�7�L��ʤ��0���jt9�*���Z�~��T�;�R`I$j�j�\UHn��jV��>ペ�J�OZ���l ���	ˡj8�jG�,�� �)����',����ϐ�t?��`��~$ڠU3_Y;V���԰P`F��K��jI��pAE�b>�p ��3Mms���5�Vs�x��@U��,w2?����gF�}׭��*�2Ƈ��!*�qqi�'>_���!�<23ß������l�u?x.�D6��W/����"��0�ޡŻ�@Q�aR�Dओ��/M�H��:#qտ�n\�#��9��|��N��Șzq�s�#��#b��z�����s܀ח�bJ������2)�esqW�.W�wU�2Y$A&%	���z��`?�j|k*���ϕ����ϡ���y��Z�������`�+!uG<r��l�l�dQ�jbW�B����ASS���K���j}�pÕ���̴�i��Mw;w�o�l�N�A=FYwxs�+\��,�.���%�D�XNp�:>�M�w�,���=��ۉ�?{�|.a�G/V�(K�[''���t��B���7�:�q��	*(��:�N�1P�ai�
���xu�"�*���=�CY�~����L�ROC^r�,r�%���N2��f�����h�Y�e��v�T���k#�w�W��#�����mY�F�^jp(L�7B��g��<Z�j������ρ��_��D������4Kdr7�<�\N�A�Pi����&�����Hx�A�g�hI�K�L�\��ӏ���P�?��E[e�A~v"�OQtbm��n�ú����{^�DŚ�B I ���ׁѤ_�դԒ2��`�X�����\�~~wo2o5}2L����_����y�[��c	�
��Z~��B����������@UbE�=���?�[��&��[P���M��&��Csǹ6���UB�:��y��91r-��$���؇��=�u��R2hZp��5��a'P�n4T�]�b3<ױ�'�XeTeZ�OP�2����\��I���$6	���0��i+��`��	�0v+�eU���NcYr��'બ�o�#�+̢���iD#C��s?��>hz�kL���&&�Q?MI�	h�1��`�n�y�X�'w���1�1�����i���(�s��/Ul�t���Ժ����*�~1�{A�0|���])��,���� ���۠ ב.�<���!<}�z�`���6���=�h@;��_�#s������~����}$�Ce
~A�_(�?�H3F�y�,p�(,��W���V�8�W'�*�V��I��.,ݗM�"��Ņ�'
$v��C��u<�sq��'p�cb�.���1S���N�n�!��u�V��=_��ŏX	�4��c�}%�� ;f0�x�p�
��e��sr9bu��Ũ{g�l�+��m׆�]Ӝ$_��Fxxs���2I`�,}�ۯ����n�Zr�ۡ�GE���!2���^���6>B���`�|��u�@���x��n�ru�}���#~��_܃�E*>`�q�R	��?�1�[uj7���t�׍^��T���ʅq��!��R���(x�5�/<K߲�J&�{�{����QNu��W���(�ѯ�~�MWc�ވ_I��yqȏ��B�kL��5&J��T��B�2_�/��9��DC���|^A1���M2���إz�>ٙ�k{�3�\�R����4%�:�::�5'^״�����]�g�`g�*��X@��G&#���N�bU(�oj�MD�ݻZ���
�bW���z����`}cڤ�bGk���͕7o����1^���1��f�(��_���y�L����na	�Na��QIP=o "v'��UZ�EbTm͓!�%�Z���v�J{�o[O����Y�&8n{fJ���ˏ�$~@Q���lD��=��,�������ϩ6 ��Ue��!L����c�x��~,e6u�Y��׶����D�=�j��Oh8:B�Nio#��7��]3x�}Z�Q�/ɩʁ/x���,Ƞ�!8Ę6}~���]�.��Y�XFٶ [��1a
}a����sY�ǌoo�FH��il.�[O���䈿��l�����h��pd���|u��g@�k��ߒ��D莑�ٹ!٪��=ԣ����F$&~,�R�ٙ���&';�[��n$������8$x�+�3F�}�yh�i�_DC{H��ԃ�s;���(��˲�G/M|�
�c .��+��Q�'�M��I�t��][��U���K��M���NR41�J������u%hC��G�]�7�Ӄ1(����j��į.�Xj��zVNh��>�/�-s���>>��E*|h$tY7���a��۫��F�MU�����[`J�#l�\��d���ҿLr+���7��C���#;3d�}Y����N�Ѣ�RxT��S��`��f�(�.�|�t�ݭ_�1>���1)�����{���VH�/O��8�SqO�|��K��G��?ŭG|H]�x����鿯���.Y�z�7dw�"��)�pZk\������m�3x�y��!��*��4Hsn���L��I�����)����bnją�o�շ��׺U���Q!��^d�v.��@�C�R���fc>�_��48�;����y�e!��Ʌ�t����-Y,R$I��GI���3���toސ����\靧D���Z��1�L�X�02ɤr/J,��5ɏ��;�5�V �cԂ�n�\�<o24�O����4��*��y���-V����M�f0�݀;E=m��1��$?ҁ�xo�[t��.�phۍ�ܔ��P��cy�n��]�@j���L�&�f��,��,��ҥ���-A��<��ᵡ(�<�!t9Ma6ߚ����e�-#j�(�	����[����(�lqsk�sz���U>�}�H��y���l�X�������@S2ֺX�����7��]h9�����X8�����R�o��_6{�<�C0����kB�-�ɉ�p��>Ze�X�K����⴦و��x/����]e��x�~���UI��Wޤ��W�L�a~���f��h���
 �B�"D٤ 2� <u���0W:ߧN"�HS �~�Z蠒ӳ����hmF�>���av�C2�z���^����1�o�Q�DQ��ed��������ڐ)J�\1��Q�u�`��jR39��͏?x$�Ց�^�����/F(���˅$�H�1BR)��嘴	,��	8�l��/{Y��$Y��zLF� 7jrЪ(����%`�`���4��?	#i��r�V�I.و�8��L�x툢v���U�~��o�V����8- �?�6v��p�Wݤ٥����b�o5� �Wl]��� Ԃ�"S�(�ʰ��x��h)S�7���8��y�'*� �1kl�vr�)6���#��Q��\XW��1��7/�r�|�+UB�Wf�67��v�׾�p=��	�0u3�,�tu@
d1H������9��.�Wt���u#rc��ޝv)�5M��n��ն��Q}��%�_VR���v.o�Kn�whB��ӹ����)����}r�$��I*��dj�bF�'K��v�(#3޶�����fd�]�OZ���,��-#�;�ud�X��B2���	Z0dts�V�́^+�%��lT�%F����`uC#_��E�T�~�4M����No{����f�OmfsY���ŷ0�ʡ�h �9��v{�7�)AT*"�G?a���l0�j�Я��XZ���_Tψ���Ca��DA|�<��6V��d��Y�t��;�̧���Ԍ������(�&��l���*[+Ǯ�=�u;�x�S�S@���.��8ѩRQ��a�8���@6$^����{��V��c�wm�8f�u�,�+pw���-�V���Lhِ�0�#a�s�x���^ٜk�$��~˴�of
�!�<��˝�DNgRS.�&sK���D�0w�`+�%_Ȍc׏O�щj�0�w�����ˣE !�1Y�^\Z��$��)�S�$и�����G���t�iO|��5 nu�1��5¨����Sx��9�* K����il�o�Jq`��D?C�L��<�x|�t�y��%P
�53�JF�һZ���>�??������ӑB���X�����4AL2Utm�CB� T��E4��i�^�(��S$b�e��o,A$=�,ne�Ե�ͪ"�;Tb���sh��*eg��sC���b�'0Fq�s˅�hU2��� ��a���|k��h��s�E��1���& C�O����!��V����6ts�"�UtO��ݢt�S\F]ژ�X�g(5_4�o��LD�rMN۝����gf��b�62�� �y������#����d�O.��0:�</�����̞�	V*�1u�V1a�c;�*./3KS�7�#���c ӵ�����캢�~�f�jz��+�����"X�	�!@����A����,1�ޠ�'Ԑ�N�ܧR|J.�]X����N���\�n֊�	9��]���� ������i���q��ho�*3`<�����A�L&ZsHѐ����)�d8K�W�5�M$�����B�䂓ɦ�;h.��so1T�z��T!ps7=<�]]�Od��G��?�@�+����4�`��/�(`�e��ضkcy�Ι��r�S�	1grƳabv��Z��?���S�&�6t�{�-�]I27�x �q�h���[�3�y�����P��>$�����ʦÛ��3y?�[�&[������6��%�La�����Q��9���So�d��A���\���	x@q�s4X�/�<�~�������^Mԥy@�E�̨ʪz���1�[#����1)�vJZ#��AEL�l�`æP˫~���H�aXS��]N�s���r��v֯��:�y�S��
u�yvhɣ���Q@���Y����)}r�59�r=�m��uk������CIBg:���m�<�
�U&�-;�)���|ZÈ�r�ms�3őق����N*�]Kn��iڈ������ƠϿ�,�O��L���Ab��:�݋7pK#xe^E\o��#r��'b^�xC+o�J����d(�����HT�x�΁��vA{�r0U,�k�ȡ7'b�C���9VG`��+ֵʏ7�� �j��
� ����z�9A��!���,��'&�m@(2YZ�q�p���6�<��>1:��=�Em-��>�2��*�踸
\2MPc"�\��q1	�����_�^_��F@�G���598��X�%�w����#��"��e]��G���O2�@�0�c���EW)&p�Bo
ݐށ��\�1�}@��u&��G�U������j~�?��-|��M4�M`�?� X��2�dJo�*���s�{�G#2����U����SH�����{�ߓ�th�Y�ɑ�u&����w'u�bVT}��D��Y_��	Y�mӔ)���!H�%�$B	M5��P	W�,�x��-�M;��W]�
O`�q�.�N��p�(k8���ǔp��� o�}LZ�x2��!�X��i~'�t*Dw��'9vW��;/]/7{�8Ixv�g\�����0їΛ�##����,R�F8��}"k��`����ɫ�q2Q�2T��ύ�1W���,�-('��r���F���I��w��;!��ˏs����4�LY�F��e4����!� ����C�w��jM���W8g��y���r.����Db�+�ܳ]y6���F�	���A�~Hi��q�*WcL��c�V�xK/���b����vӃ�v�z��Ej�Mp[����gT�����Ӣ;��R>v�9g���Ht�x�e�c_�IP6�(�f;�{8G%aW�sP������VQR�&?�{�5�$Iz
(�(= �7ύR��bz ��	@=nw��+4��^.�f�Ο���I&�Ih�0C�+�I&y�,�:+� @%Y����~��tm�u2+QH��>�4"w�0�F�n�X�a��v/g�+�Z1[<�w^;J�� �f��Dp�X0��UL�%aə0Dx�~cu⎫�=�����]�$��[��|�r��%��<������H|�j9Y��b%e1Mjݹ8a�_����n#���B����a����~���`F��WjE��o�tY���)DI�~�mH�E���F~�'֭ϑJ��fs��ߪ:�_�sD�w�G�vX�dy9�!qs��%�"{���3N���� b��$Э���l�Ֆ. �J��E�w?S�Z;�m�Q�d@�Nc�R����D��*At����������~�e�V��6����5�9�Y�	��`���Jی���"���W=�0%����
�.�`��@n��,7g 3e'R��]��y���x�\l�n.	м�2��?� ���'>��`m��&Y}3AsU�jr���<���}��&�̷:���Q���~v`�T�Mq�yK�! %�FL8Kh=�)r>p=��fG��ʑ�#���}��K��p����S\ŕ���� �F��ob����:��F�c�d��V�������[=t�uc�󬇶.^�p6ҥ��1��Gr!�3J�bs�r-�.��">&t���y/���!W��i���*���;�\F^��QNQq(�vQ����|��Ɗ- �n�GnM�d2|]Ha��(�z� �)��(j�.[e4x�Wp�S�R���2�^JK��í�J�eA��;Qi��PlQn�J�7,5 �/>������ ��:�[�O�Z������T|�y~+�x����:�ëр��5��T�]'x�NY�&���!�Q5��@�Z�a�Uc}Z�{��d�V�%�&�X����U�Ae]�kw��V���=M�i�W���{�� ������t��S�;U�.0N�:��ۖ)9�Gm�G�_՘���m�DW7J�Ѧ,z�Sl�OR�#�(.��W��q�r�$Q�y������J��f�r ��s����D�c�^�h�?�8](Y��Ҫ�0�W]/E��
�NG;���gw��񁯘�J/��#�Ng�Fh(�A��8�S��\ ?N1�^��)� &�/�kb�ƐL/x��.�X;��h�X�a�j1�M!A�r��\,X��PO�w��)�b�M?f�p��5?c���z��dK�)ɺ�p�����AH�KKB"��S���j/m�P���=ˮpNEAj��vr�p���s~X�/J��%�����$��W�C��q{l(�Z��<i�Y�;,`gW��c����^�0���f�����r�FFv��a�^�=���F�7yY= q�rm{䇂�m?c��1g��j3�
��~N幒�d�.��j�V��z?�a�߿�#�-I�S�!k]���[-to�HT	<��%4�4�M��}Q3 s����r��8�c��9��Y����� L�P�	�Z����hE�L�Tk(����'ز���l��c���qF`��6 �}?�Cɳ�%[
�:"�>sj�M�����p�&y�b�,t j��أ5H�d���멭~���H���c�S��1������*�#��|Q?�
�T*3h����r �i�D���u�%$�M�����Ф��, �2Tr�h�܎	6�̡R���Ȅ~�t�Ku2;���)t�8���(N�������@ٕB���̓�/����-<�8k2Mo{j���oH&7�q|�W��L����g��cDe��VI�#�0_�vQ�Ϩ�@�.5���ұ/�s���hf�*2y���n��Yݓa�J[&�vӑ�9�Hq캊 ��y�W�@��ex��к��t����
_� ���͌�F&w��3��je<���J��	V���⡹ç����i9��F��<0�jI�?'��������U���4
a	ay�>ҡ�q;��^��3J;��".��mD�m��� 
�wq�Я�I;�	E�G6(w=��k��C@2�Ԩ+�����r�]fn�왣;����ھ�ЃC* �2G����8I`�Sj��n�Hwpi��l�����*	�M�R}Bj=�	6u�AĐu踂�lZ�6���N��:#��U��{�#�A��1�RX����]�y�������wj�>���?��p�ҽ*������Ia�ˀA���+-�^)hI�(3å�hY��ƣ[�:�(�Y}��y�>�'ͨ�~���S_-�f|�75d�69_�������m3>͊��Ri�)�T��}�n�	���dL�ڰ�����+8��W�;��lRm�?UHi���L�u�������i:�UPy�@��b�ΰ3G����dv)>6_؎��[k���؉�ņ5��e?mJ©�_>�7��!���>�'Ĉ���x5��*�nޯ��߭	�UV�Ѻ����4����b������,x\�Ў���l2a�u����<
c��(UOX�����E�ݐ�䢲3� ��yF@��-:�2��s�weH3k��d�Wω������m��.����B��y�������������\����.K>�$"�FH�&����b(c 鑭�i�������y�i��;Q2T�I�|��>_ԓ�ݔ��L#J�c:��Kڠ33�o��4Z/�Q��!� ��!��J�u�L�Vo6֣��E���\롏Tc	X4��)�[L����f"�a<��OdJ9�!V��er]-P�n�1��z��+h(����!s�c6y�9�a˩1\4Rk&[�@���y �M�!K{��|��2`�[���E{`z����^�*j�:���*F�f��Q��X6�N5�h��Q��m.|3�T���?��צZz�ܹN6�8eO�`Dh�Gu��оzõ�%1�{�����]��F�k��(���Ǜ%5�K����Y�v&b�SlAZ�x�v�[=���_U/��>�]�e�EPq�Fa��9�g*m�Ē�Hp^t�k�4�>@*/�=�y��9lyq{-�!�3��y=mu��%T{�3Xiu�?���RJ�FQjs������@��N����h��$�����M�JaҚ
�+<d4|g�,�l�����M�F�ADBFX	Q�6����f)�e^��g$`����$ �Έ��c�)����A����-����|V`GP�]�����mYtζT�@���
��$6�I��/n�I7��� s���]y��*|����:m�{�$p��&�K5D��f�B>�f�Y��Ù����UxUɫ�`��4&�>��}�+��c2��2�����-���H4�&�!��Bz��U� ��|^\m7�Y!�]F8��x��2�C]�i?ӫ��b_�s�/48_NC(i�Z+�R�*��|�([ �rƑ����IE���P���4�0��z����i�$����,Q�K��A���pC��:�Mկ\l��w6��]����[�z�#CW��U��Π���&v�J�j��K�~���5��iv$�Q��J{2�~ՑA�@~��<@E����m��^��r��{J��34����=@^mGUn���,�x;8�03�}C�b@�o{`���*p}�8��g����w$0pRd��!A*Z�LB#�@���f�fP3�C�#�󕜩cСm�)иbA
���ѻ�Pr�g�+O����/�������|�dK�p��ߕz����(s��'���v�3~.}[�D�W`	;���UK�EpeƲ���L3qnWɋG�=~z����q�]�R��^���{��������Q��q��s�Q�TxR�	"	�օ*�I1	�W�x�ݠ�<����zH$��L�"��f�3��0�d����ݒ��f��$F������bʊ8�K"����|��@�&��j�P,>u�X�}��Ȫ�:�G�i�S��:n	���!|fA ¨(��>πj���_s���٣�������Ũ�)���G)2�{[��p�1v_��Vg�$ؘ�
U��x�����q��4�_Dh�8����n_�g*N�_�
ej��'��^���ߗ2=HwGϋJ���")d�# �^V6��#*La�v���=Q�'	)U�Lc�Y9�g���bͱ��m=�	<~<`��׉/t�=�|�uɟ�_u�?s��	����۫�	o���q�LE��?�ʼ7zɄH��~L�s�2�����;�Vm)�i]」�(�_"�BN�}�sTy���v��~Z��V]�������EwgV҂�� ,1��*'�l��ӧ���w�$'�������1��^��[xU�O�霜9�����
��<�C�;��W�JY^=����v��ok����3�O��dZ����R7�lQ0;��4�}�d%�D�7���0�P7�^��a�a�,�y�dA�ܣ���5�`?��3�/xڽ���'����mϚK͈gw�>�;��qg��"��������I�<߳<�(	��A�K��i��w���T��s��/�����ﱪ)�D͈+*�pveJ:{Z7����E�R|�x������]_�'O��A�3�S\ؗ�Dtl��}����F�ˣ�Z�@���XrQ�|��GRzD�Y��n��_9��CS& ���H�/;g���8tu#�"�Fq�]CU{�\9�̫v�L4�:�������&��^3zY�[l�|����A+K<�d\��'����"��a��/��1��]`����ˣ���u�H>��`���]<�њ>/�5�!���.�o�µ7�"���:I`����b���������6p�gvh�&_�����ԧ;WO��y���KU���3A���U�rmN�-ʃG�}5	��O����(Dh�����yE��<ϊ�}��0 ��a�wOn����:���*}䏄~�wi��3��ǸJ��>b ��N�~�%{vS�n�H����Z��H�U�MH��Q�]�m_��@X�l���J��*�<�t�l���2��4$�|vddo+uI�n��ϒ�@�p������zt���b�"��}�����o��G�ɦhfr�Ӻ�l�G�ɜ��;'�?ߧҨ	3�ڐ�#�$E��^�%4E%f��:�\5��n]T�҇�>�8�����*�/&�I��z�˙���IR��A��*����@��QdC;Ќ	�^xK�a篊L��5��Y]�JF��ެ��6@u�VȉU��ٽ�"�|�q�~�!m@�"�!b�8W�)�yNdw"������w�ܐ������A8�����Y��؁8ך�C_we���_g��"�P6�[��?[�&`_�a�@�)�F3���ލ}k�Xw����H࿗K�-��}ܺԜRQ$���{ >�/�!�V<ܚ� )�������b�\�sӼ��B��������e��C���6��� ���n�ȗ�I?�~�9fp�0G4�m�-ԻA�"��.�bc�mh��⿅;ArG�G�Xj�UFuef��6���SL{~�5"�x�$J�f/�+��̾��E�ݜ��_���P������9ND�e� ��
�[� ��do3�j��x�i q����1�B8���A�Uv�g	�3�-6�q���&4-%,��P�֐������8��?*������W���5̀�g�r��GלZ��ahT�G`)!/	&����/`��[�����=H����f���n�y��g���?!� z .0�Q���eژa2]U�N5��بJ��U̦1��e[=-��M7�ιLC/��m},K^o�r���$u+N����8V��	P;5��dNH�6�%�"s�n�Tս6g���4M}�����eZ1=��b����ވьV�ծg;�~],��ژ�(��ݻt�UwW���;~����5zy��o`|��ȫ.�d~��Դ7�GG���w��7
5er�%~��Y���7<i��)3�x�*��=����C� �5wc,�\#q}BA�p���#�����W��9Z�>��?�h���J��%-(��-�&L���%�^��@�X���W�t(2O���N��[�ܶ�<��՛���
y˹���Z�NHe����K��Hg��J�`��?������iZ+����o5�|ω�B�j�����~`���,(�6~/j�0��<�������Ψ�H�)Yh�[<}�ݜ�C	^7o�.�k6j��l˺lB�6�{Gq+H�=v!,�Y�^,�����yM�R۝��<i���P[���V�^�^��	H8�9��3��ŰC����lX	���Sd�SU�
]��qKb�:�N��I�irx�퀅������B�$l�EE�ѭ�q�\�Nh�G�8�s�����T�uѶ$=͋�%��i�:/�������%b�j.#9�o��ݴ��5��]�ֈ7�\�3m{b���*'-���s����U�k�sF�d�,�oִ��a�R2�F�!\,C�`�<�΅"�{>t1�(͇��f'���������K�S$�]�	:=���R��kTw-��/��Ʊ'%tN��&kK��Pb*=��ٙS�LP���GW:C��'�A�j���4�'Q�۝�"`ȏ�uk�J��}�
?�B&gCð||�H��~2��(�E�ԃ\��C�o"�p��SI�`��M���B�n^U�J^)��]~���)����t������]r�-�(
��lC��h�k�a��9���PB,E4-���}�3
�\�X���c$����'��vW����V��j6�*������w�Qzɱ�{�NP��u	U�dQ�wlR���jA�J����1P����Wy�Ğ
�E3�Աگ⢩�ri��}��'sk�Þn�6.�Z
����EZ��ZN��G�=�P�l/5s��J�B��!���U�lW\=��[bť��Ä�.� %΄�<4���0|^i;A� ���x���H2�w�,v>՚$�+1��A��0\��RZ�'#}��b�ӥ{"�$�K!M���tgpN�cpH��V���U�6�,�t��gyCpE�h�d�O�ց�$o&O3� \.g�����r�����;��U4��Û���㟒�Wf�l�&��eF%=/e�5�~�������Q���%`C !��vRh�>*�Ċ7*�Q"��>�����</ߵ���4n�2�P1r�Ԯ�E�(0�(�ڙo���g�U_��w���������?�@���x��H��y�m�)�K��RB ��D^��n�UA�Wh|��-Ũn��
0e�u���R����t>)|�-ùk�ߑL]��S�vߡ�{{�z�3���)��/
�*�5H����xXT=�v/ןN���⁜�
��@$}c)�!�-���  ����xzڞR�k�<�p�<G��V�S�u��3ʿ�)qc鄌�EO�E��ns&�'f�L:|��������Û��b�@��"����;\r��	�iJ<�����q�{��pץo���g����8�h��)���=}+'�w�"S
b�C��5���h8<Pc˂4�Jf��v�:�L��7�NQ��7;��=^8�߲��g=.��Qt�I)�:Ԋf"K)Bi����)���$���B��8`'Mfݫ4T�9�, �>}���Sq�2hNB����jj�`�V����U81h#c�B��������HT9�`��D�Fx�Ծ�T��6�{�=�Hę0���t\�d�{��K�4+A���,�-�޷�<�Q�0p��p1�=@��+�;H�2�Ʋ��p�y�����p���&?�'�SR�2OQ�g���{Z��%(�Yb�9f˾3�ɒ:�X�.����,YdIo���N�`�U��ۆ�� ƤNz�q{{��*=�"&�����{b� ���h���f��i�5�ϥgw����na+�v��^c��.�9���=����,��)���"���a�Y-s6��r���H�	E�	4�a���+˩_v�	�K�_�*�ͳG��@V����#�BL ���4��$;���*~�!2���.���$[Ԭ��(�*����)ؙ4(B���~�#F* T��6��q@�QO_>�w�/;nD-��Q �r���Lb����yA��i�R�Y��}Y�Ӱ%�E�p'2 '��K�D(՛b���DG��
���B1J�؅��3wL��^��L�f�n�.�鶴�������IdGs��Ϛg�E�|����1�m3c~��d�ff�ҧ�\T��!Q����.L�Th��z�p��_ 

+uN���%˼M� s�S� �rQ�D{��Ĕ��લ��/�u�����'	����߲{џ�e�ݬ�[sH��1Q�R<����:ɻ�'Z�К\�0�@�$��U�z�~2U��m�C���:�bf)E
���^�g�hm7}����A�LK���n�^U��c���w�6������]�j��ڋԘ�@��E���f ��i�Џk@~'h)�l#�)��D}m�t��w1
W�Ӫ\v������§��<�
��������㨋����<KBOP� ��?:��Դ�hg呰 �+�����t`�]H'7��+i�}�M����JjJ���`.�r�k-���!>�P�y�针�0��2˅@OBӡNw�?'b`n�#U^V�VRC3�C@̎%�=��t�-�������`�D�p�_��=���������k�D. > ���������պj�1��/���^��U�['������0������;N�b1�m-�))�vL����"yKZ~�uvXp��iM�%F�y��\��x����&��p�%KY|�{&���v|ߊ�[��\ȟ���_?�B�0�&בFBd�Q@�8�E����5�#�6�}�E�m�2�i&�_��ז=z<)�,�����gUpr2��kS\�oQ��jg(6ݫ�<p�	�52 ���;b���T����Kq~Qh������y����ڷ+l��E��\K%:A�����\,O	��X�@9�����x�M}S��1�����8�2\�.��'��)WmTm��MW ���DA�bm���x��`a!��8��]N�at�~�0�sk�,[�ݙ*y�s����j�r-+%J ����!e�ޅx?�rBN��Իگ��.B�I� z}gQ4�	��G9��vӎ����ҬB�b~��\=�	;��4x� �%��ѯ��q�����S��0Y�#_>�w���ɾ�2kA��]J��N�u]'��+��[= �p"�m`�>��z���̨PO��&i���"�jE��~���DS/G'i���OxSޢM'��N#�T��U-N�`��m�GV#Z��X��*g"�W�/6����6X�vwZ[<$i߶�[W�(s;�F8���S{��u�@@�/Li3s�5�D=��E
K�o�ђ�G�=�N���U��yҮ9��%Ij+שa3L2i	��~f�&✝���;��B�z��f~;���>�*��ҽp2Q��s�G�D���CoLm�yP�L$��b7��i!oz�SX�����$��쏾��A9�i�#"�B���<N���E�/�!q�]豾�IN�V�u�r=���}����c���LoPd�X=���P$�8,?_~n
jo��p�ޠ��tAT�_���8Y.�^���U��j�4�yZ�����]fΒ��2�!�UJ=��"�a\�!럤�]�N�5
�cvs:����8�P������S�4��Qh��CǍ+�aMܥ;��I9@*Z�p���j2F����5�n���2��O>P�vl��Vʔ}����t�ܜy�(^1�xY"���HM����Φ���\h�ZV�'_�:0U�yq���3�������*	�hE�/��	O�UI�m0��d���p�X���#@t���zH�*,yy���c�X$��0��M��d}�^��A��|���8CIP=����h{F�՗������mM���Ƙ���_mj�]�r���Lܼ�".�e�Z�x���`���d�՛�qpĳ=�X �Q��uL�P0�X��p&�w �E!Ss}R߬�MSw�`W.x�J�]�Z��!M�^�F���"�����b~g]LC�5 �u��a��ۧ���BU��eཐ_I��R��<�6p�1?��j�Y�������w�z�'v�,��WYl�'�֫R����d({��e���gxV2�v�-8;7ڍcAT�FG'�`w�CՄl�l�]��YЂ�h��Wm���Sψ1�#$=2敉T]kI�soC�{@�]��������IL��I��c")�,H\���q�#ҿ*鮩Źh�H�w�O6�ˌ5��R�����rkV�b�-�����h��6�S�}/�\}�w&vuH{�5�f'D�P�����Q p\;�	B�My�gl,EK�%`,��$�u��`jB��r[��V"�;>�_e�EA=*nP��#�������	��� *|(�R�Q�Y������1����K�@��ѽ��|Ue>:�'��"���;�[���ɺ���犵ڝ�e9�c��
�DN�tƇ���2����v`M��D�)�x���i�n�TJ����sx�� i!��f�W�@�)�<�n���Nh���-s��s�����mX��^z���_�2�03h�h�� 	�B�-{��W�Ke�1v���ݫg��.��{���_��d�h����5{ Һ�P'��+(����Қi��Bb�I�FpɪBrr�#�W��?'�V����x/�����ڤ�M�9�Z�I!�f��Q�ŒA^�#4oV8d���wԚ7�;p0t?�Hp6���B%Ya��m`�[�7f���:�vq��u�@)U�1C�ruAx���$�o�=8�֗��)�5�H�p���Ni�&�����5wJhݫO�,?�;ce���Qm�}����]��Ϩ3��|_�#н9�5:��/���כn�U_���X��9&Yr�;q
"O^���Ω�3q�êZy:�%�)�;�<cl�M�6�C����m6�_?n����u�]�x��wW�D0���!�-��.-M�c�yzn�̅�i^��N���c���]��6�8�N�E���G�L�y�mΊ�܂���;Sΐ��
O:�D���ر����Bxyt5�5�<z�A����~9sD��\D���e�=R�-�3SxG��@20��gɑ����0�Y=���-���>g'[��C;6�rZ�e�*�K��<�/�1t%��]^n�%=U�i���@aY����.�:�	���7��A4H~xU�3�7���hM�C�X������1���)9���⡦@�1禯!F�z�)6�?O��Y;Z}��Gߠ��0J�+�r�*��ms�{�
��*�X�g/��UɈg��\�P���i]�ٚ�[�V���,L(�\���
���gm:�k�8'R�#!	�ZI�Oe,~z7)��F��� �Q2��7
|xhŇ
k[���F�
v��m�U���.PA�l%�q�F�{�1�H�g�v�H����� �{�>�;&�p�XS��z��R�!w�t��M�wN�&b��{�Y�� ����_�!,C����ُ�vIYR#:�Kw�i���^ڟ.�1v�6�FQ&[�4+��B�idɺ��aeV�E�`�����k�_*l��A����w%�^�WY�}غXcF�qy3�yA��`����urI� o����V4����E�3������Q�MQ�/����7�ZSmU��;Cr�*���rX�p�
g@Ƣ*dF��yc�4=Q����曃?�rob)�G��=�R���W��@W��s�V��9�%���F6Ǖ�(��tV���徬��'��I%U!��`�,m����E�糟>Ug7Q��\�bD�8�ŷD^D(�U�[�ř
����5����`��R�-�	��Qzt�c`M�\����+��O��|�Wp�W��$�Ru�`op��w�Dv�_}����KF��V�c�r�U�u|��~���j.��8�h�q�J�F�L��钼^ �	&2�Ӳ���b̶Ӝ6@�uLW�Hh��jA����U��S��9�3r�
�O����m��n���-���Z[�8��X4��U����uX�[���,S}�Ų���)��y�'"8����� ��U�N����������E
�t������3TD��6�h8���23FHu�߶6�^;+��ÍR'H�jl��x��>���;֯%�L9-7����g�	l�5d���ݠ��!�t�X���g�k�ۺI�bĸE���KG�(�{(mk�i�ev�2:͹�~�.-ɲ��C�Q��Ϧ� ������� �
[@x��h�����U����e�5'<�g�q��1S-r2��iz���3��t��ֲ�%�f��a�yo߅���.��&�x(��-�9��3�EV-i��A�XD���G4�yO_)�j��P��6�ڵ�QYD��4^ڃ���L�=f�QI˗9O���A�{b�l�i�xҳQ��1�`���~c�t���o>Q�YXa&���£���r%��!
U�N2�(��x�9|Sb����XD��㙂��D��5�H{V�{��w#$X��ɍ��L���E�"�H]3�=#N1ID���3H�}�|;�z2P+;vlAs	�K�����:3z�1���c��;��k�1�ڃk�C;�n��4K�*6��!�}SP�!q*_D�E@V��w���:�p�B�����fSh����Q�2f�����g��x��%�"Ν-�Ȇ�w�#Q�ǩ ��{����Oa�ɔ�8��bn�Ȫ�_ ��� y�K�+��]��L���#��ٲ=%Ɗ��{��A���)ĲxW���-��K!̛�{��K����t"�F~�z�p��O�G�&7OLy�$Y�/��ey0�����$���e��)���I|�_�{��=���:B:q+՚[�駋�.2Ih`o�b�IV�'�e*�$�,Y�u���aW��R	���W���ũ�l̶9X�&<����Mg��T~�gf.��r�w�5( �a�ƨc�ylk�\�q�f=՚��7�\[F*欞WR-~!RbR�u����/��	�Y�!eY�1	�t���A���[3���J�7���~̓�B��d^�[^��o :吖�{�%�$�3�r�'��(��F�h�לՌr�/�$�Lw'-���a�;���vH&%-����n?�sS�+��\[,��9{z�� ����ȩX�.��}�j���$N��U
Q����tk=�D�?������Va	,nP��^}���f��:J_{�P��"���\	��T�q����]V>n�A3`�q��@�+}��̉��fS9�9�43=�JԈ��B�%�X�e��h�f�2 �4�jL�0zO�G�oC�!|7�IV�!}(kY'���Na-�����:�p�֤>��#���/�-Щ�AC�[	���i6o�@�s�M�(���>'�k��B���X	i��e�;�ք+n^��i1I���< �����a�A]��r���0Z$}�"\��O�.�q͂������$@�s�`�a��(��.��!p����@	��0����{����i��'��=�SJ�»(�%":>r�GB��<��9�6��iK>vZV��������i�7���W���*�ʕ�)ʊDW,g�R���Ȭió~����;��@X�-:�I��_YTXR�s����Y�Vho(�4�a��+GrXp�K-�[�b��x|"�%�|��z`58��ZJ���'���� �/[�B�|[me��I=L�#�Q�>���L�v�f|��F�"�V��,��\h���L�$^�7��ޮJ,��z��MV��W��F&����m(��)�O�=s�G�t7��gP��^YA���ԩ�����"'�T���*���=2p�������}"��e!�����X�Z��e���{E���*\WE��=j��-\HKcRhL
G%��.�$h,��QU�H�aʽ�*����V��$1���8��e;��k&fq޹x�T�8
̅`D��BWl�"��i�T�KA�F{̎���I�����������S�s2���O�� ꇲ���B��y�'-+2rD�h��GVKv����D4m'�铕�&Y=7=f+��+����y%��q�=�~z�sw�~y/F���\%<Pt��=�ֶ2$va�0 ?�%����٦U��y���V��}���ί�(ve�y�ߡ%zk�����@%Ia����iJ3�M��EzSٻGG�^7i�f��w����)�T�`G�@rV�v	חB<V̆�\���ŝ��EDɟ�3���w�G���u`��J2�Xw-��"B��p?�Sc΢�)�2q�s�5��AH�`�P�^dh��%XP�M�hG�57Զ�����n��o��?�h������f�1�y� m����_�Y_����eO>�
u\�[�{�)��)���z�i&=�r9���t�`6�a?��p����`
�[l�LzuR9X�Y���UP������Eh��L̺t��!�j�����G���:�R�j?�}x*���4a����+�?����FJЪ>��\4���)�c{�߲�rU�X�;��&,�[���bu��7 ͟�޾}�*��6Ǚ��P�}»5�e��]�ƹ�捸�D�~ڻ��Y/���Hl��9������+�������P)c��9F��ج�k�Չ°��s墷FN/,�"=�2���p��rI%cȔ aA�	T��};��l{	����暍I�RHd��>9�AB�T�0�t�:wa1sk������"Y�Z���e�N������#�W1�"���:�W�E���}��&�x�3e��t=>��Cǜ��o��̝��"j~R��w�$��6���g,,�K,� �U�\a�t��]����3�~X�O-=l2؝���m^� }��%zÄ�2��5��#���1�Qx��� f��F�e^����h�\��!�qiְ��/����2�ܵ��2��ƁI�0�7F���j���q(D�I��p"�
zl����_�_�I]!��
�������/��������vJi����]u�ЃB+�}*W
ݘ3?�������܍�ŏ�ʄ%��2�կ	�$�pM�t��-��������g�'�m
�}"�` �8��!1�7ԔA���C��@��<��I�H������Xb��V����Y�}�����9
�r]����=���^\^ˢ�j�F�Z�H��~3�Z8{�E3 �0)�9>�� {֒��@�kŏ�#goj�ůC	�^�0�c���s��ܗ_?`	�����Մ*��13Ϫq���й���)�3 חy��k�Dv�Zl��ϔ(�G�XK��Ĺk=�'�qg6MX��*]yӉ����:4�;py�x����fOd[ؠz��u��p��T��w3�,�|���ծ��Y�S���E����/��qr�.��hgzcv����W^���d���!o�Ɓ4#Z9�k�&8�'��s��H���g�?�ؓ�9N(��B�b0[C�K�ZD�'{^a��_�>�\�.]���-/+�U��m�bl��yh1Ug4��?�y���M��n����BC%3�@�8}����#v{����V�@��?�����]�P��P�s�	�6�Y��+%�x����\��3S�l�p�F��;�FY\b�K��y��*�깡�F���fz��}A�����[�NH��Ê�{���	H��w�*#@�6{n��ѱ7���� �[{��*�ð�l����t��	���c�V����ӊ�^�I^�QW�l���J9QyJ��F�wXr1*5�*h�!��<ѩ�Rdi/�R˗���$z=9F(.��<�	��	ժ���xM��G8��8-�
�	i�[��j_����� ����mfT�)	o�D�N�[��X�q�}2^��[y�!Sck��i������|�h.����PJ�܂r�f���)�T@t�W)�8Z11~I���P}o��Lqݞ�f����:��N|��K���q�n��bG��n�̬#���|܄ k�`��q�D`V�#�C�`�"��G$�3���Z_�"�����$�.7�䫆�1
�,/�<��FN��������1�	�G�Z���i�Ȇ�ؼ�W�1���\�����@�i�>9n�l�.���:�jӒR��|EA9�H�C<~ْ|��9���m�
OƘMg2�L���ur��o��S��Q�+C�������{��늰oVe�=�����t��������F�23;�K��=[{�C�`:���֍^?l˙G�h~е�b�%X����k�ee��_�)a*#Y���v �*�Jۭ�nG%�M`��Xd�c�*ϊ�r���,A�� ���)Ǉ��\쨒X������O�%�<D3�TEC�֗B�Kn���f�q�zv9��h�O�BŔc���s��G؅��ZW�a�rx�>Ԛ��|��$%� .��{{Aq�a�8�5�-�B�3�	�p:v`��V$���u�d5�v�Wf�'].2�]��C�C.:� ��	����cd��x�6OO&$�k�Z���}��[tj�I�i����.�͑;y|'����'~bo��}m��k��p�ˆ�O���|¡�������̧ͨ�.�v'���T�N��Tk!�O�3o�4�R[a������(;�k(>�(�h.�~��s �XI���}�����wܫ�m)��(7��_RTM;�I�!E`�2�#��wF@��G��|:���ea���%�e�O�5Ј=R_"<L��!(\�Z:��#"K�
�`J��M��Y�h�M�J��	8}W���f�p�tX��^���|����4�2�_�h�� (��?�#p�.Z�UI�_7��(����jy�6�!��
��{?zDG�����jzAے���B[���$��t�]��-��w؊)�^�u�m/7�+�Y�x���%v��h�6��C{̬! �cƥ��i���\�����f�dE��<�e���J��̻j"���J���X�r�3꫋���z�b�Eٴ~뺢�v�]�vw�N�	���$���v.��L�+�Q;��7�2)�K����������Y�s�I?sEx!(�\�.^i�u���8M<�R�����(�⦚L��Y2��=���/t���$Խ����N��KW�5�7U�]�n��c�Hf�i�y�"K���a�4M�9⛙���ӘD��{޹�}oV�M�Qg��8B�6 
���#��m=g�ç�w��o6^I�a����.K.�D>9ȡ�*��`��vꧮ4YC�wcd���y1���~�q%��^����0�EfY�+�U7�iy�b'������BHE
����}�>,�\�8��N܄G�UdAo�y͠����q�5�Z�3�A:t�v��е"�Br�y�������_R���O?#�x��=AqI�p�dOYE��N%�?֏V~,�ǭ���j����^[�A��Z�UZaڞ@�a����7�%NR����5��H�I-�@�z�7�-�!s�P�Tm�Q@��~s��
G.�l]V�=�\�ïZ�x(U}w �~M��=��1��ኂ}C;a%�M���F�Be;���9*[� �^�B�3blmW�\��:�����S9���E�~���r��ð�C��K�g^T��X��<�X�-l-Mץ�ЂZ�B}~'�:����w̉�,![���w�_4s����lIq݀��^[kJ3M=�8�W��5A^Vg��Y����^P� �D#�pib��i����̳��Ql�ڭ��9F�`N���~����#�QOwm�_(W#�,�4]���V��dT�@<��l3�?W��?W�w7��ۀ��@�W���SqK, `y�Ͱ&O
��X�D���y���6��h��Fel�L<T�YI������y����Et�$ ���smݧ��&e��kv	�k�U��ůz%�IX��D٢��$�|�H�\5@���� o,������w���,�w�/܉TL�F3�$�r�H��gu�%
��N���4�p����.���V*/����sJ�;��2��I��l��V&�I����,Yp;�DKv�y^U�B�M�Z���y������T�V�e�����g�J��~�
���t�oj���:�q3LL��y?x_�]&oJ��z�E�hķ��<�M��_	H��W�o���
\�T]) � #��Gv�s:l�V�$�֙�T��EދvkT����(5��I,�G���c_J�o)q7���~�7��]+r�9���~G+J�~q������>��F������j��F�[�K��T�4/p�* Z#�a����`s�?��Kt#N�%��\>nw�Q`p#^� ��	��d:B��v���F�s�@��3+�s�v��a&$)n�lj-<K��<���xMES/�c��X�2���`
�B�a��(|�Z+V�9���[�`ׇ5Ÿ5�j��0��֟W� T�C��o�=V�]��s�@V�����
T	G���7�Gb>< �~��`oyT�L�b���!C5W����CX)��9 l�@��)5�� ���m������9����pcͼ�T17�B2f��ٵ;}?s���7��,Il�T@�9���U�Ӧt�a�З��(��g�!8�6�^��:R����k�}vW'�*b^;4�- ˤuZ/�V_��� �1RF��Y,���V���|��S�
�Dwh�rv$���r�=֓�c���t��';��S�Zp7x+�m��V� �3�^4H}a�H��w`(>� m�U��4��]���� ��SJ6���/��oȴL;�.3��P��+�UR�1��F6��g�oc��oWࠩ� ���n��S�]�;�j�P���FK�7]��L ��FfJXD��5��l+5����\韹J���r��T6FC�EXt﫮R}d��O����xk��A>�����.�7 ��S���?#&r-�!L<G[��{b�IB��@��n$d��JH;εm�n�[,��C��t���.�ȭ��zw�<����S�L�R8���p��(m��h�����kҶq��~�.6YԢ�kX�d��[��4URR��a�;-�DSΐ��r�d(�o��.�<<�PqH澇Ӟ/,���I�)
uWe���O����9W�4k�wV��z`m� /f\�g��lS�}HwV~���.�#��:�g�\���9��'�ڣ�DOɻ�b3+�&���ɟ$6x �c��;dPy-v�G�w�twN-�=���X�`w`Z�(];(t̞b{�I�U�D��v��>�0/��j������ľc�?&�4��0��A�dVQ�j��[��Æ~XKP ��<ND�ҭ8O\"��p?�����J�2H\���01�:�X^���t�*"�;�sf�����Mצ�G���k'�ݲ`�#���~��(�|�7�9��u��8��9�ᾖV7����NK{�%�ij������'[t����������~�{Br6̳Q!��]����	��,	�Xjn,Z|�����%�U�6�o���g�")��*���d���3���qY�2��刐��	�2>��<v�蠚��V��K�zi��(��Ե�I�#� �$��LT�d6,am��Uo6 �A�r���B���ڞ��@�p$d��V�]�@����6a����|�i�)n3v�v����i���l�����SXngXX>W� o}�ƪ�0t5�]_��q�S�Y��-�ho��ܩ�:�tv����+�Qz�D����Q.55�5ߥ��d��������Z�U��C��}މ�"�V�c��TS1#�n5�w+CK���H��4sS�7ݯ�>�u
��Ջ��SË߯|9�Oӗ�sa����9��?7�MY~��l]�Q�2���Ї��t���!C2v`����"���%�m�h~+�ṧH�j�D��*����&a��.�6c���#������ ��M����&6J�����$~�o�r4����$��#�h���) Y���k�������<)�E�.�-@��w�k�<�$$�ٖmȰ�$��	�����
�P�ѱ*D�G���j�A^�{쌙�����9��u1+r�b������~2���u��c��1�`�V`��χid����-�2�jL �ۘy?�ʿ��Yћ�AK�dh���)G���y��l����s�D����@��d�*��B�+��%�u$��"�w��em�B��(�l���J�% \�7*�	��
���M��`�,à�p���m#�G5��P����)�}#q�~3�G���	���̧��2E��&�)���L�h�r����:��:ұ�)e�{`;�˾�����*���o~r��(�y���ӯ��S�x��}�t��'�Y�v��ڰp��8����{�� ��a���B�}��C�*�T�1�p�f��k�M�P)U��s�@G�+f��cS�8+���@�BV��j�\>SQԘK�4�xK_��b<>î���MJm��Dc�|���>r�GU��_���#`��F�L���W�gVУ�Y)����*��ĘE�����o��4	�R�SMLW�0vQ� ��	8�J3��l 2�Ņ��e/+F�3D8�Έ����q�]��b�����nn%�V�|A��!�' ^N���sc�3���z-7yZ��ے�k�;��g���o0���l�G�y��VCQ��NO�Mޛ*|��!J�Vܥ�f�&D�V[����q�#���N���df@�Ie��:�8��I0e9�v�)4̛1[/�s(hS}r���p� d��e��>oXu�B�Յ�@ٌ����� j���l�԰j�	9�sJ>X�Zb�]�.�'���!F����=�&��Fk [yP��M�
���6�g��(���蜍:�{T��Y���\�� ��U�f���=����6�"��A�_Y��[�����q樂�%�PX�T�vq��3���;�n����F�=q�[j����u�e��1U)��:I�A��G֒ԓa"��	��Q��<)���#����c*�.~��g�~�q��Z�����U`
�jN�o<޶� �7-����&�F�>?�L��X����Z�,d �8���5%]�64�;:w����"�כ�<r�Ԁ�(�d���3LIZ�}6Ua���^�B#Lp�zܛ�,6o���=��`�U49#�a�[�({���f����n:D��4"R���$ۋ`o��XkO)��r`�2��|���V {T��e���+A��A�d�]Raף��`�=�{��0.-Էɓ��*�	a>�w���_�ln���_������@ٟAꬱ��\���m��
L�'�Q3��5hR�>�mh��B�G����ߎ�]X6�"�o��@��\�%�O	xQ^�Wз����0�bF��@��xCn��@��#t6�I����<J��5н��d�=�z���1�� A&��_ZC������*貥����w��pL�},I�<�脗�,a��0[VCS�����w�`
��>�b��f猒#���G��85^�7D�+������h�A!b81�s��l�!�c��;T�������iV�J�㜵��B&!Y���R�S/$��d�2�]9��x�&������藥��h�v�!|!]��44y/���O<7ѝANM�-͏�-^J�)�{=`���3R���6#�I����^�:p��WRc��!�?�$(X�o��Qx_h�P%r0�O`�]YrĨ|��Y��VO|}�2U���<5O�)}nn����3(ةJ��c�Qp �m`��Р-)��T�K�KbOW	0��*vC6�g�S�M�{dS �D��&!1�W++}9���2��Y��_����. �m�T��BLz;��f��݂�v{hCV�t򃭵Z����#��7$ȍ\HS7�\����4w�i2�����ӝ�z���|d�+��,�5���%<��t��G3�Ij��zlu���s��I�sru�a�)�1|�V�o�ǹ��9�v-Y�TK�k�,K�=��lQܔޙ<��OT�A����J��k��n3|��+y=u�����Z��欐�B���z獝t�A$�
���ĕ�3�{�%nMf>+�;�N�Q~��:���ΕTWY5TRf\��_�ɪCiyC��j�fp��P���%}��uj�Ck������9�⫑a��S�\�vTқc0$Ҥ�P����p�󺭅�0�@N)�lx~� N�i��e��pusey�{�����76����v}��tXa29�קKZ�F�^�TT-�&l٢Yg�({i�H�{�è%p�f�D��xF��}_-sx�����0�4U�N�
�K=Q���|����ьp�dD�d�6EH
�<�!ޠ�7��$".��ә���+Z�Y���xG�� ���rI/�?Rvl�!j�TJ����ֶ�'�k��+�~��<�vA����}`C�Z=��G���/�A3��JL��}����UV�Gk����h@gpxp�y�Rա�5;Uۨd�Q�\��ޅ����Mfr,z�l�/y^�>�����M-#s}-�j��R���KEd���vl��K�EU_�66J8n"w�0����~5���p�2��+ц���hX.sg���������r.�+ǃ�#98Fl�@�{��<�0S�j��x���B�f���TPRL�uQp�	�z���k��p<�7�K湢L�ƥ`���N3�,��2u�����i�WC�.-�����)�|�[$��q���;K�:+ˋ�� �k�e�z�����q]@� ��NA��Ti���{Z7�p�[��v9�ݖhk\�%y���2wC�aȇ�Ll�u\f�����'.��¸A);`��jn���Qٳ�_� A��ν��%��%D����싁q�t�4*8��f��� �WTl
� �`"��9�񮞯�6�(�&�$nE�40� `�e4�J�t@�wP":�j-��p���D�Xؽ^�1��B��SݣK�v��^-�l�v��.M~��Kgcz���<� 1w��F�2��v��ZpKi�˺c��%�g 0����ҟI`B��t�S2󿤂됭�G�Y�w�M�҂���J������ž$K�� mA����f�Ps��Ig͵�Ϝ�������v4���g�y7'����Cy�"'+��o$W/@���g�&3ڠ'W5�m�w�J<!�ť�y�~�7.���\�s$��nv����~SA��3�Kp�I��N#���'��AwRV�=n��m-cƢ��f�$j$����Kg ��x�"���_�E�3��AɰV��l��T<]��hK&��)�f�{j�6m[F�����0�,��G�a*8���BT��<N�Xirg�2�V���W�-�;�x�s�o�U�� �؁�Y���̅?�M �q
;V7~'���	�q�Fcj�J���S-�/=è�K�FW�}{�,�!�؎���`��m�CK�376�i9��b�M�b2��Q���ϒVW��g�������	�L��מP���׮�"j��E�܀�%4�K4ldW�O�[�TjOp.�jz�1ߥ�0#�%�h{�GS�}h�IX<�s�=�_���2�h�g��hS��>2�I��QסX @n��u�r��1Ϝ�Bu©��80&��8��E��c
�x鿎&������8_I��L rx �XA�Q�������X1�d�9i�:�RI�O�Bl;�s��45Ji40+! _yJR�D�N�_*W*C�C��i�V6��>��	�L*��8�8�+<	J0%:�K:ׅ��;��W�]�D�k�a���� d�c�ظ%�xǢ!-^uy���к�:x�b���i��ki�B�%�9���\9%��X�>o��Q�����4�/H�m�sӤ*+,�W C��`��p�����K��e[�q�RH�S�r�xG��6 i�@ �t߈菢:�����0ma0��n���̔�_�|,��q�74������]�`a��2���ت�*#����e������+ƶ)W&�Z���l�f���1�,ǟR,���B_>��g&9�I8�#�Ay��%�|�C!� � �FQh����'n��_�YhHZ���eJZ�gˢ���Y���sq����SU ma@�����yo'wXM$���:]�� ���q����@���$f��d��#��Jƫ�|��1��k�Dܺ�C����`T���$A��,�HE���<�=ML�<w��	>�r�F�&���n�;���@V�V�~[�Wk��T}=2�o�˓[%�w�4h
�w��nR˚<O!�V9��-�۴��+Y�OeO&��/��{�*$Ew$����e�Y�������a-'%����?��s0b�z�^�%�.0��-qU���dL��	0���&n<�?�#Y��_�t�z��lV�?�>{6�#!�n~�ܙ5aSHZMv�B�l�n��:�T���hV9O��=Y5_6��I�]ҋ�!����2�@*���2UG�x��p�dY�[orP�z��i�Ul�͋���׊��w�D1(�'������szW0׹������p5�:| [ԕv����
:S���A��zL&�"B�������b!OF�3anu9�c��J8(��{I�]T\�QYG>�;f���0 ��Z%|�e0��M��������O-�Rh�������/oC���#�x"o�<���ccO�k#V�b6���\�M�?��SŎ��Hd��3L�KO�ƕ��~�w1�x�	(DҾ���P�$9��2�(Dj ��C읃���4�]�/�A�hti���t�e�S��o��oi�yя�JWFw���4+��Y\x$�o�B�(�p�Q/�;:�����f��]2yx|82vc�Ѕ�����d�9�0F��[��]��G�@`�U��b�߈%,s^��.#>�����s���YnX��LZ�lwV�G9��JŹ]�]�(V�%�ƤǥЏ�F_qA�s}W/ý[=�(��<����W������s"F@�T�RM�K�	�yI��<��&��G{�=�t������o�H��ڍ�
������< ��Z��EOa�w��.�PB�j�Yve�Vx�p��S]�;B7Vt�9b�_����q�|7�:L��7,zA�H�<pv+0
_�m*��<,m�0�g�NE<��3��L��:r�:h�w��mb�1l����{�}󄻍Ga�ڕ.��.���a���Bf�>���6>$eJc�{�.b���f�j��SSe�z��nh�6s�����[��-R���?:hd��qK/�dr�}�$�H��h��q�4�� a�n��b��I�!Y���x�4u���a���X -h8��R9��/�e���aM?<����>�!��Y�������)B�n���W$�T��i3���0���z��XeSa/�Jp�
���E6��J�Mqk_��V1L�d�����!�i۳"Z�����r���:���pL��ֹΑ+}���W�'�5h������+žZ `�t�dy,���/�� M�f���niK.��4���ŦXwI �%WP�\(TϨ偡j��KK�BG��z���/M,�]g����x�O=B��OH+��`�w>IC�f�X��5 ]t�a�R��6��ځ�vKm�@5ͲI6�FP� �{�m+��*���|�/$$��D��hGF}���[M�I���{�)����Ξ��5���$��\YU�h��
�J��c�l���ʏ^���x���ώ�0�`�3>2fpN�&'�4��x���S�~�7�s'�tJ�ީbF��Og���j��F���>�4~�ϐ�}��8T�Ӂ�l��r�����:ء/L�*���Qf�%� ����eV�߭� ��+��S���GO�#�	�uف�?Z�������Zو���V����s�9�d�C�>����.���MK�S��늌(�}�OR����m����Ze����ė�/�]H�u�[T���4\�o�&��K��#�xvʸ�n���j�w�r�P@�q��S�a�y~F{xN�~ǭ�m�������h��b�m ���O�-�/^]��G��ǹ�Ωs��'�EBy��W�L�u�����Axʌ��}��X�w��T)k�ɦ߄L6��qO�*���y}A��E<�/����1�$SV:�1g��m-��Z��Y�v�����=PY�[�@|T�B� ?Wಌpk{+��I������|�λQk��{�)I��`�Y�t�4��{,�17�l ,��� ��lv ����"P�C���t�\rs{�l��:�v��f���-qߝ�����J�>�m�n{�=[.����b�a4U@��Hf'�".���(�\�L+W��96;Tw�؛�ӯ	�f�h�#)J�b�87M����׏I���¾l^�9��'n�坹?���q�xRViQ�i8jM�;���2}�o�V3�@���,�>ص��i����`�j5��a~m�ѬρBƼ�����"�a��g鵸ei{�oo�R#�/��j���t	[� R~���'\�nכ-�y�/���T��~��l���0.�v���i�f�%�-�2�c�!��q?���ь3l�f�(GZ��00����@��'����.�g߮����w��3N5l��)*2�aSp�3� �6�{�4b:[%F�t3��L�
���U��x��'���v҇>c��;Gt5�R���^ƃ�̭r�� b��_���$ޱw������6p�����?X��-Lt�ҕ��A�[��G�D��o��'͗vdX�6)�{N��*�65k�\��|����]�ٰ����;�}/rŏG������HUX�$��13>�W��P�hT!h�g T9a3佻5��8����$ݟ��I(�1��.X�ZR��y���v�,n�k��v<�	B�w�{u3���f'dA�*��V�������������+�`�!%�1�<&�K��N��񊁜@����r������hS=5K���L��E��Wx�C�2qRjv�����
G�YL���T�_os��*�� �C�̽1�) k�k�b�VN���LB��[����!ĥ2�|��<e�*E�7}�re%�ph�W��uӬ�����l��|��XD+�g?E���64��i����܋"#����՚=w]�x<�=7]��.t䧻��K"
ɛ�}kj'�фhx��e����1�����n�hbI}����2� �D�Q�XJ�A�q�ɔA���M��V<e|�#b��þI����Ǿ�傎��ϕԽh��ě����6��u�!�2�t���i��<���,��cZ:��֪�Q�40?���A��T����^J߶��yC�6Fz�2�;¿�Z!�%D���nn*��e/#0l~̽t�+K�1'���R���S(�PI�^�K�/'\��I3n�N(��#����/�C�;�����0�]+��:�����'�{L��K�P��s�kVLܨ��l�l�[�Ci- X��R7��-}�����'߄�<��h�?�T�q	u	M�Dr5��^�w��M� �������;q�;ś������cٽ7RʩF����*�1���.����o���ߵl�@a��zX�^=J^�wri��X�!x��K%�A�� p�D�>0-a�2���0�<�m��B<��=Li��H�qkb^I=&g��W�D�u�]�U�H�e���Ť;m�B��[,�����6*]6B\��D	(�aQ��r����w1Aj5�%'�t�U�0�����?l1=��t�}RL.T��6�3[]�O�UBcT�|�u��T	\7���9?�>�o��)��XEz��'��/\뎾��L�$���a�+��:3�R��xօ�K�p��ņ���E�2������- ϼ�����L��绅h	�Q���2M��l1D�{���h���6�1/S={��k��!.	����*����J4Ӑ/9�8p�Sr*ęy�c=���5_( �杴@*�4�?����e�w��t��jװ{e�]� ^�K��J�J� ޓ�UN�G�3O���j��̡��)s�/g�}^���YR/>�A8=��'�$+��A�����n@ܛ��Nvx�K�+���v�.�_]B���p z�W~a��)�g�#��f��G{�p &/��Ñ�Tl��y����R����H�qߡ]1	�SV��s��p)��dU(g���}B@�gl�4���;�=���2����J�^���Q$ϔg��(Du�l5�2f�[�|��4���3�L�O��.�Խ��"��C� � ���B~:��@c�v����c\��;Ur3L�YU��M��[��H��:�'�`U�Y�ϝC�Jk�E�Pd� dz��b3�^���Dr��sP�@r�[{��Β1��@-7�X%�t�斝���6�vOM2����(�J��-dDwL�y�^���J�z�#��:��S���3B}�>�/+��lE��}��M�M�Hح}��݇F~�s"o�}]�BL`�ػ�Uş�����-��'�[�B(1�;�Cq�
���z�0<h��G{D{S�~��1�>��B�ޯ$�����SG��>q����K{ae��5A����8�L�>p�k�����yVO�V��N��V���Äu�z�f�����f+��t :��	�X�9�D%�Z!<��"��Y]4�\Q/��~��`[��ҺR�ݽy�Hч��2��Ϊ�,�wV6c2Bs�i�w�Y�?v|C�v�$Qu�n��jE�S��N�\�a͟��O�\&�jBg���S��x��r9]�D[^�{8Y"�]�:�QsvӈH��vEE�����(���.��8�|��3�kC܁"Ij�4.YY,�)q�=�c&�^1rw������1{�9���)b�l���ٯe�jW��ə�<��XvH���d7kvJ~�y�;x�?"�u��Ս[a�Y��.�U&��h�3f2�@R���U/�����ݤ4����ʃQ���3lw��R�;�VB���C<���R8�����W1r���`mZ�Q�d��E���,v�u���5˄���W:I��������~��[M��D�Q���&k���h���_�rH���H�ыM��7���ˀ���*?뾪{�؟���aG�ܹ���u"�\1���������R���;�xB���>���`���\QU�j	-j�(3t��`"Yۛ�ƫ�W+�Mt��FqgҦ����EO�Q�~�5H�BQ)Q@S�42�e�UA������������
��,��М�OEM;|2��)r���SA{�������`���M!Q����svw���jؠ�-B�V�v�|	����� &:��K�^�>�y���v�i���k���9)��!w]Ա��X�~.�,����"`��"yb�#|����/L�}��O�v��YeR���.�#$LC
8A�7��QS;�q���5�¦}S	����4sa��7�I�\}�����
�d�w.bG][��A�� �F;��vE,<@IM������e��B�;(<���|�1��5����ϔ������p��''S�%U�n�g��ӫ��'m2�W�63}<�X��Ol��*>Ml�:ƻ�$�)oVl9=��ƛ�'Y
W�i�*;������S����#)���\�C�i��V���BɲY�>u��S�.��b���<�K������=9۞�S+6���+L[i!�5�RX��
����iCO�S4�%�LC}Z=�a�.�Jx���!S@ !�������?�_d]���\�.ᚺ���\�`mk��ȉ�k�4v��U9�A�c��&iɅ�(a\��I�sP� 	�δ�0�
s>&�� �>���U� p�˼h�r?�p�aF��C�Zn�[�Q27�CҘ��$Щ@(�}z�����b�|��7�[�w��n�J
���H�x?nCD8���TZ���@ ս`���bH�h�!"~���|kJ&�&�����ٕ߻�y`B@������x0��w��3�1�¶Ip�665�Uc���9���3������mp)����A?eX�u��#�ܽ��0��ių��h-\�Yh�nuư%��a��Ă�0s;����^G�)�;�/7�#�?��9�O����_���/��T�~3o�l�]���t����I��r!y�8l�v���6+�3���AW'B�^�>��u$wEM���ǾD"�#�.��G�y�P���	G��;O+�����L��<^�*Wpj�R��jf|�C��_���g(��<��8�9�zY�ɴ>��e���o�wDmB�QH�磱�}>1���(��y�d��p���xD=�(�X���h�<�q��S��L����Ҕ��;{��߳S�91���]�9�rv"Z�?K�#^���8�.S��?{�@��r�����ȣ��哴������p�bM�"���f�6k��{�FxTf(}�Lw5�V���;����W�C&�CUo��.��Ͷ@��$l��� R$��泣V�/|fy�\�X�~�l�����rbɕ
~����͝~)p�Gҍ�.�7P��0x%���~X�iJ�^��EW��8����m��Q����?LtG����L~�鋮!EC��X/��֩���w8G	|�N��oA_��I�H�'�!����fҮ<���,�Q����-�u�Qm ԙJNRm�{2�g]��h>�`�Ӊ � .s�ܭ��<?N���T�v��Yq䬐�Ɩ��=7��w�۝CF\%�x�	3�1ѐ����[�y��բ�:�u�Og�&��>XU/x
ŐrGӌ3��r�tRS��f�������ʟ͝r&��[X)3�sP~�2S�u�;�o��<@��S��şx95�Ƥ^;����:�`��S�*̓�7@4�����G���yOUf�O��L�����R6��Mؒ_{@T�?NAg�j��د��&�D�\�rT��x�(�O��i5�A����th/Vo��2w䭃:�"�h؋3��7;2y����F!��v�q���铯x�irueم+�q-0�@$�?�R��_�z�����T%^����R)�۝3��M! b�Ng��a`��W8��⾻m:�8�6t�P"7��V]������5�D�����F����@�x��zU��6rk%��fRh�m�vS�)$ݘv ڃ5#�}Ж\"����)݈!	_�����L"��GkzLY�gI��Q�F�&�e�ȏ4�g���n\�N�����b��1y���N�K.-ŏY�PM�4��Z؇c)��6.��v\��L	�;9�q;G�4K\� N%�y��X*5Z@��c�)0�H�� �PP����)�d�q�aG�[�YB6���<��u!���ķ�J�a�ʹn6�Ta뇡:w�<C�	p�>&5��
1��`�m��c&�]J�@+)��"<?H�k����Y�xXu/��6�?R-��O>�U���͓����a#hu
���'�7.���(���P���-�۹��qж��2=*k���-���</�f}�>G��	C��TXWf%Ű�>{�����ʢm؅u���(��W5Q-8�o�\���V�H?(H-�@�<HwI:�&�����CW��	F�R��޷��u9�Ց�=/��ۍ�O˕XGg�� �`��v�CS�F?�{�P)`gs����1W����cǨڏ^�M���X�����Ƿ� �	�A�'�ʘ�*/�ZbN��-}g�m�|]vnm�C��x�ރ��oCI[���ì���#Xɦ��i��{E��	�<��B����,Ú(Մΰ�_�VyQ��f���7I��L䨗��l;D����$��AS��������w��N�����L��h�ȁW����F�$):�lU�An8�O�J+�1h}�}(v��f^����A�χ��0#�=ΛξD��*��S�&��܊D�`@*$���NĽ�թ�H�,+N1/�CE�
������`o����_��;�Ą����%��a;wҀ��:�]M���Z#��������p9��]X�mk�~	�|M���Y��`�"�c^;26f)ӹ B��6֕0L��'�e�9Dg>����z��_c��8]���TS�L�݊�-1�]�)lL�q�i���
��[:�������cՠ�U�|������la�O*YF��?�vC�	`>�6=#�zAF�={�{�W9F����-�����V8���?����O/G
�-"�B���&��j�
W�[�?��u�\�q�n�|~���r"Sz�N�~^i�=y�J	~��,��]����~(7�U6�+���VJ���0iA2��G�?��#�tlտf�Y�m��m�"�\��M���Rs���<̝�P/�����Js�����m4���"Zg��Q�{�t�fr�Ƚ��z�>�t��������4����J�:zo��7���.iת����U<Oӈ�Q�%�Eĵd~��w^��z�$�ՐQ��}�f��_H�h��ǘ!A�3��T�*���a�LTQ��%�F ��R1~��,P�R�.�D��	�|{���h-�(dw�{������--0�P��5SJV��s��}A�T��Lo,�y�_��G~/h��o�+�0~YP�4S��b������"�>VhZ$��DN�_��EͶ�f�#ȉ�Bǳ�P�ǖIP?�M�+o]Jb����`��T��oW��<5>hʎ_~*�l���V�����A�PAI3���ߘF�E��3*	BXi-��{���`ߙ�b^zsr�ܽ�F�s]i;J}����#9
�I4��@��88��Qrw�Ί��\������3��ժ�]���953�C_�(��>|�"��exmB�Eq���(�����vQ���QC�Â��6kM�Kg�[J�)����|^�Jx�1����B���Q3��OR��6O�8ӝ�&�(-sP���yƴ
<Y�7߼FxhP(�R`���tw'�_�ta)y�5�853!�� �*�K�֪�/��wyW��6Q�i�.�D����N�u��U/M ���:��C���.�<͛o*��ۗ<��Zi[�q�;.9Q��#Z���a��j�"����0�H

���s��	b�"H�B9�2'܊WR�=�M_̘O�!/�WS�f��
���V�kU�|��NsL���O֒Z�'fe`���|����D�u�y`�$�v >���"8����-���*�zc��V��� H
nb�]�^}�G���y�3���S ,�;eJU�X�����⽏Kn\�P�E��YP&l�9aR�'x�����V��%|4�����W~)�y8�н�57k\��)8�:��va��ARz��<^K��n��&��=K;�@7!�J�+�"ș�.!�F��,ӯ��F�M��%wem��L�c��e�uܣ�\���V
�iH�Q@: u�T�h��/��<&5�����P@�䵧��mI{��:sn�J%�_f�dNt�ϋ�8@��j�u?�t�)挾���x}��s_@��������B����K�nB-ڦ:L5z��oF���@��f᏶�M��p�lԢ9S�.�U��0Fq�U'�:v��@D1��X��������_�T�1
�HB
��i3�K�6������2~?(�H����Ӳ�
cZRsI�m	�Z�x�p���kʇ%D�|�u�h���q�BN�2h�<B4h<��"��w�]^�[�v���:�]-�&"�;���,��&���n�|�-lSL�Y��5h^K�$:c'�Ҿ� �{�Hu2bd|�}��f�\p�E{��~��� :��1O
��r}\aHw�ǀ��"O�$����}Y˔ܵ��$,�m[�	A�fL��N�����u����� 4�
��B8_��낢Lt�X A�:/P,M��*
�b��ʮ/�T�E�Q��g��M��DM;�9�a˙J2.��๨�ɶ���-���I
���2�~Y��[���lK��V�{t��al�q?:�I'ǉ�-7r�w�A�R4+O��	�6���Ru����0v���Q#5|b�b��N�CZ��\�9�U��1/Ya�o;�J#KG�=���cB\oj^"x���>m3m3����@��l\�J�(�ȘV����Swby7�g���B�g���c��lHm�U��*3��fyV.{ma�_/
����a.�;?�.�� �y�e:W�C;'�N����P:b�3lm�LP
*�r�ԅj���M�i@c�Ψ>�P�P��5��h�r����60V3b����LV��'Kbp�%hiO�PH~_Tvh�+�XM�������	N��S=���j��j;ݒFr�dіO)&�5��$�@C��fY�[���s�́:�7�kV�_�ӯb�&��<�?��_H60A�Q�jJ�1wcO�IJ���*�)NG�ZIzͿ�D"��a������*Ԡ���@�h����Xt��F@�/i��C<��}��!�ϓ<���KGq>ذ�u����a��8#}Ҿ�@p�'�1���Q!�t����h:�*�j�ö����s�ÄW�m��:�GҾ��7�p���LC��@X6?����d> ��B{��؄��-ش�{)���r�AY%>,�r"D�AG���n�Ĳ�(�C�xz��h!}�#�i��vDJ.��1��p|�#`�Lq���&��K��OTs��}���G�̅����O}#�?��M��
2bUK5����[��Ҷ��\�X���#k3w��{�����8��&�������f��d%���T(��ݛ�TY�������B����HJ���֜�EȺ�����K�SRX�$@����x�X���o��T��d[֑�SM�_?����a�������L;9ޞ7y�jݰ�7�0y�ݡ'?�=�J��+��ː4'�x}�T	��<B�{�I��7p���2>N}#Qd&m��˯��{u=$�j�ޙ���>�x+G"Xd���C��1�PXe�^P$�#�u�#�jzU��(���w�S Q���`E�Jb]���0��R������[���-�i��LI���w�˒� �C���f<8b��z�9ѥ���}��Km��/�ʎM�
MOڛ�N�`QmUz1'��}d���D��*Q�U=Hk�tb�AWC��	R�Q}u ��� nR�<m�.n.m׺'���ۘ�E� ��.����tO���Vmܚ-�F�!+��Y�#�Fa�2�-���՘*H�e��,@
�>��XR�d���zf��'��I�1G�ˊ"���=�����M9y)�$>
5�ev��(@�/$�U��j$��3#�_UW��U%�E�����ݙ-*��Eg�Q��'Iq��,�P^(N�dJ�� ��s��m����>�����&RǏJ�fGB܏��/ ��1D�#���^:�Ğ(X�.d���ȝ��<(t�m��fB�u[�o�^�e$��9�.4a�'��fz' 8VĔ�^�8���	M�F?�ĕ�����x��J@�X~�C?R	�y�3���0�3s�ٕ�֍q�j�K�<6�ر-�(%����Jiˌ�0�N��8��ҩy����OH���芽����K@�j�.���,������d����7���F?�a�qr�{x?��Ɯ�����a��\ h �b,��i�`�PCZL2&�O���MT��%�*F�����_kVC��V���9h���zqר�Ӏ,��x�%-�rO#CZ�邟6�*^��.��u��B��S^t�'�0�d�\�tZWs����Wx�Sa�~C0�&l"7ۥFv3YR���db���(�8Y����1����b���|qKƐ��Nl���M&��
O�XCpM�ҢK�ս*��fKΚ]��Tr���\�0��^M�0�F\��dh���a�%�
�ݛ�w�%�����L�Fd��t��CO�Cr,cµ�6Ǉ>����	2��1�Շm-�?�}����Ҝ9z�F줩Wfi�]��m����g��(����%J�SBf@"x����8�AkY�ㅺ\7�m�F!m��K-����͇�1�p���	�<t�����^��Y"�@i��`V0X9�����uCX `"�y�U�B��LJ�v�����+���m��Ɓw�������VP�d��& Lܟ'��|��J�H���V�i#Щ�tx���
ce��Y����/p@R�;����c�=�qYe�}������}�8b&�\�����ك~����c���G{g��+�f�Ht�e.C�7�̯_
~e�ޚ�����l�a9��=�bz�0��AÐ��V�K?��ܻ�@�N���mW"�p��~�wJ��|��{�����z�}���!�=3Dth����!��<��°ĪѭG���Q�Զ��(4�&g��������U��-Yn�6���m�u_}���G�*0n;O�7��m� (k�D���S�Q+J�3�Ew�w0�V���Jc�\莿4o�	��D��d���NI�䧷?���R$hff�C)7B]��h��,��e>�5*��|BnҊ��s���]�9z����8���CG�"2�V���<Ԓ�6��g&Qh���+����T�D)y�h!u+�qJ)6X_��>D.�\��ƂnM5�CU�ey
m�� �ӍU)�P�Z���%�R��\fAhpf�]1%Vk�Q��}$� s�~g�	����
�m1O���y�VNz���LY�`ވk��f\{��^Ym-oaǛN��Ʂ=��Ó�[�cf��(���|�Ne��Ec��Q
����2H��}�毸�a�\e 8�-�7�H�]��>Wb7�����UFE��:qV���e����ε�Yzy�~�;]����1�H�Q�h��6����ZrUc�="5R�b�׵��Bv��(�rU_F���0�����?��5 .f��g��C�pS�Ƭ��x�e\�aP���+M�����P�6)r�p���D���?��N�����E���.Mi�!��ȗ�~}���Q�����<�h�'yM3�������H0�yW0'B���3-d���5���٬�@O�6���LL@ӻ�F_oh��*�A�P�2� +�?*zǓ$z}Y����c���Jj�T�oǼ�1�B�����<1�@�켎���G��r*��ߴт)���(L�V��Aĳƻ�8("����ƭ��iY�R�ݴܠVB��F׆�Vx�1tnF��{����p����U��8����c�ӏlidL7���M�
�YOK(��=2��
��l6����-R ���a�X=J��1���í%��#4�^�d �	�҉�=�|���vf��S�9��)��IS��&k4����QR�\K��M�: DG�N�"�o���J3�	,�f�eˬ�EK��Ȫ�=�Hu�s���*4%�9ٰ�o� �k�Br�o4�k%�kA�9�c�\α'�E�B�G �% ;m����m�������C)]ZL��R��v�O�
��CX������O#��]�Gq�f�q�����"��Z~x����vVn4�/��w綍(v`���D�^Pm��Ok��ԕ8�^�]�T�e$���GO <����p��oWhۑ�n.ٺռp��'CDci����I!���b�W���O��;'�����Q�ixO��\&��;v�z�QF`))N滗�N���R9��*˦[���L�R3`k����I5J��oHm���t�px�bJsC��I
G.A��q�b��5|[�1nh�m{}͢����-�t����J�J�(Z<(�9�ۣ$3�Ã8�8g�s�D�� ����/��5[�<"�le^��7+)ug� 뷠�I?4 }ېlU�唗|�&��&'+̇�g=	���"�������~�n�%U�������V-ؔ�"��M�|��X�f�`+�%�>xWӌxB�?����L������´�1�Y0�5ÈI]�*N_To��������Q��͋kI����jo�R^� ��vT���7�=�ZK�wl̼�����䉾��&D�6�G/��fr���Y�n⼘�s��u4���O��O�*���F�-���%�!���I�?,�0�h��V��wSh���#�uD�S���V驷 u .�:Vn��Ɉ=1&�� ���[�F�<�4ǱD��Мة����!�=)]�@[LWy�63.Q���}�BO� ) ǰ�q}��4��c r��9�e�~T䇖R�����U髙����.�X�_V��@�`�j�N�a��F5G�6��T4��[�ql�B���-��Kv�	�3�98ܰ<�8\�c',1"HJiJE4q?�=���=���ִ���L |r2��&�4�T�≸� ��~>��}�@ONڹ~�G���q��M1p»f���Ti95�� ����q����o�~������7����l��t5^ -8$��D��9�Q�6��/z��P�ΝD������>G��9�K@��aSIw,|x�!m�?��ֈp7��H�_F��!��G2J�o��xQ�w�\3R��8���y|k(jُ��+�L��i���.B�16�j�x�<��m�ҝ�=��e@K����8��_4�����	�a���E��ԄX��aQ%�^i9[r!Pk�)8r.Gu�xu��jRف0�k��V��΂�\�]f����f�Bs�O5`�&����&K������ՒU��?�|��H���I��Z��.+tv	ڬ��mt��7)|{���f��y�2#S1�8�����A ὓm0���^X������-:��	I��x��"K�ѓ�A>P2�ů4}֒��#e��C%a�i;"�Ԁ�/A�o�.8���&:�D~�b�s�W/�[<���g�_�2z��A0�P�h2�]i�����f�����RW�p��
3baqDə/ͮ�]�T��(y�n�.������y�л��5����T�t�����z���jw���­ Q9�ЏE�#��� ���	��%�F^kf�GI�R�N�Fny_$�$j�d��V��f�w��O>D�H�8�w�R`_�[�z'�M�-��;�l
b�Ԯ+J&�v�3@�-��|3rF��T 6�BW^d�u0���}h���&D�\�&
g

A������I�W�ډ�t��hWM�I�)\��<�ڃC���O2��/ÔO*r7���&/]�z&���m�\���x{���+2�{LhXȻ�Q¹�O}���{����%u�MLdB�Z��T�W�P<J�e`��p�]x@��k|P1.�w��b�"��>�Ž�"H8C�G�#5Ac.��Y*R{��KɈ1e?���L��#��S����~�����۫�gBa���g�1Xq���E���@�7ԫIÌ1R��\x���5���r r�ja��3�����<hk��W�;��?��J���m�|I�Ⱦ!T�ĩZ6'�!ʷ"0����X�by��{���ry+��	���>ް���}|M.z���Cy͛��A��:r��u(
c�!'Zo�X
����#�Թ���*펦\V1���+v��y(�>&�����^&샐���F�T<��:x�2��P���z��]��Y#����)�T}��r���@Ձ�G��
��{nX�kG�����~`�U�B�C���0�x��ٜ�u�%k7Ւh��С����Ӗ�s��b�����o"�����98�UP^��V��^�(�%�4b=���7_�w����zꆌ�o���/����?����}C6lOI���y�7ֶFiק��N��*@���6��b�S�A3*ta���<�6ۈ%�H��}��
��,  Y�P��fF]G�� ׌����x(Aͫqιr�땘�w��.RU��$�����&"�g�X��߮X���(��|��F�.���1dY��¾q�]j���;0���n�!wX�
D�:�����4�:�	��$���,�����.J��}-�XSQ k��E�	.�k�c
�ln&m�`�G���H`�ٝ:��!�`�@��y���\S�M���W���D�Y��]���c�+(SmX5�n���ڏ�6����*؆b!36$Ơ	�aX���_���Q�-]���BG0��A?��66�7I��N+M���&
�N���<��k���"�9K��S1���U�;t�։�z�ҿ4{��;0y����g��3kIT��W��v�B���E��q�x�Y�
�E"r�����8���c%y*}H�_ ��Tb��qT�L*w�B݀�q��<6�7�%d`�x]�%B���䯞�Y#��u�6ǪPQ���h�&��\=bߊ�: Ktj9�ATn������)��~�[�L-<�J��XR
^���W���(���?>�r�Y�`���Zԗѡ���R����;�eL7�V4u+�c "e����$6�!��8�^����?F�C&�f�'u"8SČר�N�p�6M�2a�&��4Ȝ���	�{��UO�څ���݃ۺM}��c���g��S����i4�����{��n�w(D8HΓ-QZ<^�����[�1%8q��/bJ$y|��Z?�݅q��;�̓�v�� }�ׅ������,���)܌o�h�w�#�KU�#y8�B�6�ޅ�GZ���̽�=O���U��	�&���.�A>�K<�9Ά>�1��fo�b ���qr�����W��� ������Ab��]w��B�!�ض��3�Q��)�f��!a���q�=1�IV
J�9��[��܊�S�ʌ�(�iL���	�Ti�ImY��H�s.a<�@���ًGL_��m!��;�ּ
���mi�O�K�ū�����2�����Dꨖ+�'�%�C�̉��0��� irO���lmsvx�x'D|ې9�?��n����$�(�� ߉�9T
�,T�W�h����N����Ν�iwNd�S��-_��(�x�u�P|$��Hu�![��ש�y��J�T�a�U�p*3�Ķ�"1ur椚��O`�� h�I� �ة!������mTi��"�6�+���F��i�?�Tx]��HF�������Ы��9�-���Ш�\e�� V5�ുM m���Ųb���w����",g�L6��ˇ�\��DY����Rb8�V n������K�O�Q%O$V�����i}E=��=��.LN��e�T���}�FC�g�9p[n�#�T`��XP�> �X��2��7/ʬ��ղ��E�����l~�vQT8Yr��@o9��n��%�(1�`�c~�G���/�����n��]�f��
%Xb�\�Io���m�Rp� ����79���F���1� #��ko ����r�G��7
]��v�$0��W�?Ҹ�R!�>è��d�˓�mC��BvNtO�MKc�?dOS���x��M��o	靖|h^�A7Mp�����@{��U��%�'M�ܯh��
'1�t;­���uy���鳫.V�A�4�>�؄0��fa�ܓ�鿦8�[?��j���e�� ����P���H���Ҹ,�
ˆG�a�?t�*_� �W{YS#h;��#��RZ�"X&�8�-3��|��m�bP�A:ؤ�*�.�B����L�	�վ���EF�i,�!�:�t�[���5B� ���K�Rg5n��.���LJsE���;[Vϳ���=cZ��M�u������c6���������"�����m��oA�B�e��5����'�!	���'/j7�x�{�9�Ex�!늊$<w�� �=��=��}e�'M<݌��$1�	��Ī���A�ח��E���u<��y�^���j���V�\n�4��P���s]��K���D�u�����1��v�4�<�J�A|��h'0���=����`���&j-���.A�GeڤYQ�pq9 �)�]�MM>Q�d���r$�8[O��Pr5�p	�T��NI_�a_e��0�:�ZJs��,�L�2>{G��}WI�B�^>�0N��s{f��W�L�
�r0�ME��fz���&B�km�K�U?�����0Ǖ�J�����1X��U���wa������m���>���퇦�Ԯ
6�$큾��E�� �ʉEa��n(�f��F@Ed�ĸ7�^uO�D�+�S4��0VBFx����3�ϝ���^ʅ���J��+:�(�}�r��D�ׅ�輇�<�橣����E 9�����9���D§bVǓ��]kr��>�P�H���M)r��Y��%��f��p��Ϟ�U��F���9n_���Z%��n��u掤���0J�?i�!��̳�̭d$�zp�y�)���[!��ʟ���c)��r~|��{)��i^�g7= �C"R{��,)^��y�`J/����b_��ה�>�ǘʩ�&��<�FA`���ڡJ��n�F���i�dx�-����s�����B&F��
5�t �g��� H6k�j�4��p���;ش��z�l��v���=��
�Pe��g�l��Q2�.�_L�]��}&�}$�߇��׷RX�|ȓ��I���l��ƣ�˿������FEfs�o���x�~��\ ��&_V�o<��s��@*��|cm�!w��XMg㿒�����i�"��8A��i��,��[�5oN���s�cD<J��C�'���.�{�S�|Jk��K>Q�3� ��L��D��L
�}��r��Gp����'S�iŻ�a|͍[�n��N���+v3�{��h��=s��Y��|S��cԉXT�������&����\J)�Ԟk�	Q<��&��H����։���v,ϵO{�mT�Lu7ƞ��^鎛=�U��	��c�9�u[T�ϱw��_�!gT�d6}���69�2����y\��ތ[#��cP9+c����$��_��P�gl3��$]�\�{%�#c�҄���%?��F!��d���A͋�4���B�m�(j��U:��`�Cԟm������J���d�ETSѩ�^�lAݗ�/���7������@&<�O����"��o�"�_i�:�lu�i+���	�2�g(��)���"��ck
�G����Bj�#��5k����O
�Y�͎aL;e7yz�;���9���١��O3����y�o��yU��Q������תJǞq��mf�h�i�4�΃C����cɢΝ`���*s@^�c%��x A��4(9\�<Q�����@��bWic��ż�j���;�ۇ�f�+J!���9K����
 'T���;ya��!�5p��n��x%i��������'�%9zU��]�bVs
V�_�)�"Y��;�PQRڢ�K��A�=K�� ����[؋{"�r��X��X�
��<p�q�mv�Ƥ�h���n��f��a������?��|����آ�*W���6��������F����DY���2���"�z�}�*3���n��rg�0�M"��~8�Z47��{e	� v���x�8ۅ���p�:�I�������3����ܙL�>=���v�ry.m�zs��-�X%��v�`Ux�v�F	�ڢ�1�H���1����z�h�����1�x�VH��*����tl����^��m�	���La͞������ݺ�04�X�����Ԯ6�h��`d[ ����!>L���gU��獧��]3g���Y�̻e���O��{s@�]���5�^pL�`0��rT|��F���M(���'J��{�߶�L�6�����8S���'�lb4R��I>H^���T���9*� 
���!�/g?��@�Z���p;i�/�v2��&`��i\���d
�E�9߫������%@[�G���D�
�����8�K׈c���¤�^ݳ3�$غB���D�����(rE�`�������Ϩ�oM%C��P��`�Q��Vj-�s�O|(7w�+���+��^r8��]�IU6s�r���
q�=M��Ǻ�낾A���%v��3�n@J��ӑ�?�]$�)��vV���('�r���n�O��qdګ���J��~"�K:����+�O+o�
����Z���4�RR��;^��UX���.f�=lz�Aڮ���gЭ�n]{x�Ҕ�HBc�/'-mV�`�05+_��CV�?!��ׇp8�Oj߃#]3&����Y��
j�|�e���HצX�Tn�v�L6�/As�� ��`�G�sQ�f���a�Ϛ�?i�cE�3{��b���t�������g�1�뻶�$q�S��+�+�t���%S��
[�A��5v\F~�͵�]7�\�	U�Тh����R�#�o�G�w=X@2��"U��E�a�AL��8�u;7y���^�~��c����A����ZD�`W��{���V[%#Ճ���s�?8߼��V�"����-����D-��<�Y���@fΧ;��da���&?L�ƀq=B��rk�tX���U�R�;^�"q8���ʖԁXg�鞙���4�t�bݦ蟧���_}���,#�4��х���@��Q.�64:R"�K��u,��a�lV�c��d2�Mc�Ԑ�k� �f0�W�@`]���b�	����pj��#L,;��7"���Sȁ˭�4VU��Z�)lշ���T�"Q1?g��z��$:�_���cFVǼ���yH\����P�޹x�f��i}�}C��I0�ʝ�<�ǀ���1X��ؕ�}�����т+yb���@�H����?��?o���zi�ǒ^��R�Z�S���A�A4D��|���s�\�9VV�n"e$Y�Q� ���
?ԴL��t�2�BY,�)D$��g�\ ���ʧӒ%�c��ЖiM Z-������J{w}�����'�TӚ!KL���{V4�F�����)s��j��E����Es��*�ESǹr��i3 ���(|��B.�0t��>L�~a�ꋈ�>C�$ܔ������)t�=�"v���&KU���v��ձ��f�� ���Ѫ�u��Z?9�M�S{�	�6�6�Dꥸ>�����j9y�@ݓ�6��d�tȸ"�]�����e��s��9$dE�
|Ĉ��i�`)��a�:��EC�+W.:��`1�*H8�mk7���i��6�+�U�:�+[[>ƟŞŦ��]�䴙��.�+��M�5伢{�z���!H�&1�YX��׷�	���2'8�ؙ��L2x���Z�=��T7�j�4�JZ)	iq����l
!\M)-��m�&�$�s��X�(k#y�=�&S�	`PA�r�d�i�rox,�i+��pP�.�&�F�,lZV�wkO� �Hte65�bA(�t������
O��0����p��s�h�!�["Z�2���2�pMQ1��yU��i
,�!9���qj:��8e!� �C�cQ(  ��n"��r�b��2��90�S������a;�m6hZ�v��5	V�D��ʏ�ʖ`�q,x{z'k`nk���>yWs�#F����t�[�����j��1�@����	���H�I1T*Y���QJ�WH/��ڳ�o�6&Ma^�mX�/ h�l��;+��m~�	^>F�$}h�x������!�3���p$-
}�*�rE���k���,)چOlҲo"���F����P/�ѓ0�DV�	��cNX�⒗����qX�V_(�d�����(�@�p]�:�]�cN���O�,����:�8#����,Qً<������U���As���888d�a��T��P2�ʢ��x�!4��h��8�Ƨҳb��O��ї2��4�u�)���������d��~���A����RP���s֜����� ݻK�U?����=�}�b�J1&�����Z��׮tL����su�0>�*Ak-�?{�j�ND��9�j��ZO6km�\�|�(�0�e�-#鈈���i�ֹF�ȭ��K ���7-�^}�T�}2��R<Ω�K���Gר�+�l_��c�*�����4���ٲ�Ex��Pj�Ļ@�z����H��$�
o�ށ�y4��(�RO�Y���Ѷ~���wx�Y8�0ы��B���m��z����z���G��V�������4MǑ%L���#铈���)k}��1��
�M��8��6~Ug��"S�n�e�Ϳw5 N��t��q�/A67q�F�?gG����l�k<��%�"��ԭ�)񗷟������gN��p���;�9�1%8<��&s٢��;�s�h䧌׹0?��v�Hr��^���T��?�L|�ȊI+I�����l,�2[Du�a;vSh���[!�b�����}�g��1�T=�h�r?^'�?S��b(�ċ}�E�=Ё� �ƤVL�.����=�Q1~����?:g� |��:MP��J��ά1^=�ʜc`��:tzЇ�iNP��J������S�F �L��b��q7�V����a	������4�S�	�?OI?W���M���`��1�������'����-)[m�^��B�p\JX5�f1�=r�|Z	p�%��n~��>�쬁����	�b� �?�W@��/����TB �h���>��j &Ƌ��#������e� gQe��x;��� c����O1�)�8jW�'�K��3�6O�u�3·���g�[EE|���I��7��m�ן���}s��zo��kR�yՄd1��D���ۏ���� �y�:�BP�)d�mH�g?�l�vl����=�eZy��`du+���\�u�~�d���葬���5�c[��p���֥݃ɻk��x����`c���zo~�£B���������F�r�鋥���W����z�O��׼$�� ��	��fo�l#3�#K�]�I-�(ќ�#˜�9�p�ٱ>�o�HOQ��^쀺:��Θ_ԃ.A哙v�&���	*nAbwK�˜:|'���B�_.� '�E�q�_�.GW�5��ꋠ뱽+�'��z�b�H��-Cè��f��.��;!h�]�j7������`#���Y���9Q�#�Q�v�K�!-
�\�?9��g�m���؄�b����1!n*/�-�<�ا>7h+��٢3����f�cl�UB���ܗ.E��V�����I�X���B���^(,�쾲]��ǔ�(EPc��u�)�\d�(lCE\v��`��3A��tz"�*+��`2����-(D�N��[I<$�?���~�=��o�ݻ�u�	yI	�D��C|�׏D���-���!QWwz)��\ê�Q�u�ք��	�]ҝ#8E��C%��<}A/R�������U�z���PR�y+l����V��%��1Z/FJ�1�ݶ�;^j�s�uf�����߀^���E/z��c^І�� QG�,�?&��FF���)֓�<�|
6V�$�K��Y���V��(�ͺ{z��d� NS�~��ϾHJX:������C�c�cpѭ��[I�&�cW{ofZ��'�1p�8K�Po��ʎH��5-��r��`��"��#]_c��-4��<�VJ�e��<7׬;E����8�|`+���'�{`f)�.�z�B;��⋈'6J�u?�t��=d�� ������p�R!���.9G^�; ���f�HY��%N15�ʧ}��l�Z�v�{�z-Z����Ȁ���՝�޷a:�������Y�r�QY�ħ��a/�b>�u��Wo	ҭ�<Bux�~�n(�b�4�/�j��� 7�5!�U袄oȉ���v�QHPf��OI��Jw�Q�y=u^�.lF��8\� 6$�֟��>��>ұ��n$ǯ�t��H�X8������C%��e)��}V��n�z ��y�gQ�
CQ�RI�c��xg�nς9�u���e}�7�����s�V�=��ק������M�+ȍԔ�=��aC�C�ɦ/��uy|�smO���B�3�M&���kr;=��N���@,9`��|p�Wa�Ez[p�$+�#�G�R�X�:��T��Qg���[s2��^�Wi�ۯX�8<g7���7�ڢ[�����X|�\��b�Ђ�P���s@��_0Z�e\�u�����P\V���P7�#�[:��EA��肣�u��}o"���^�͌�����ذ��&����<�y@��4��ڞ��bA}[AM�'x$SEp�H,���U�j�" ��VgTuW�c��kA���Q�����/����#gb�{����������Y�!%��R������?i������ǘ�)���� t���=Ci����N@�*�K�?��VR<���7I,f\im{��_­�3�ܛ���M��l����5�<���Isc�s� p\;%��s�ą�,<�;X/���h���3�]�R��9,��D�-�2.���o�Wr��գ&�e�{�i�Zp����'M";:�	�N��2�vPF�R1����6=b���� 9��I+�ڡ���Z��:�0��&��5LFfr�p	�a*J�݈��j�Q~R��ϔv�$�M��F!����3�C����z�'@#^(��g5�{=S��ui������xh��zu�/;3�[�0�&oW�}��M:����������MJ�t
��!��<L�A�C�|B�����lBhN?��:P�~",e��ђI�:������Ow/��)	<z����=��FYe:!�K��i�ڋ>��Ń�'"��)��Je�*�ix����6W\��T�o�nhJ�;��Y���1�;}լ�����x4RSW6���	�9)y����	�� V���+�!�K��KJۨ��R8�bQ��>�$�>c|�Q�Y��`]`��8qj�gc�?BE;��nU�uU\�|Ð��q�~����������t2���L����������B���t��3&�:Ei���W��A�09���_�m�5���a�х�����9�GJ6�.�T���"q�T:�%�����܁{�$Q��� b���ogp±�Y��E�h�36-�t�=�� �Pw����	�h��l�Y}�:�ҙ�n�*��������L��zG���� �~.��z]�~S)��/=������Mc�3o���8 c������3��� l��)6���?� 1<�r�a*����Zb�N�i/��F�,RWx�_���'��df���y����#sM�dk�o�)T�2]U-�b*�iy� �{�Kk�;W!l$�ڦ"eG�ap6��C��]�A�1�ŀ�䋪8�#�uш�G�$�Y�;�>[	�OZ��.�E�Zx���>,a�%4j/ފj5�$�pB���|��钿�69*�"{Β����a����;j(ɷ��9�?ק��3�{-*���"τ�F�Q��cWf�ZB��{>�����5�>���Bm��E�����
,5�����Ľ�Pr�wD���,�Wt���2l$�>����P0t!����$�j��DB�5h� -en�;��tN���N��Z;�Am&�V�؏�6b�����2=�2�D��&��/$��۞x�]�~%�R���� �W껡k�����i��{�;�V���;�;c��f���i"U
d�&�nڼ='��7;�gs$��*�Kw̭.�7���iIw�H'8��@��L�T�"5���8J<sצ�и�?N�Ib���kR����.Zn�yj��X_lH�l�3�Y�C�O��4I���8���S3���!���B��_�L�5����Z�ܪ���2쟏+@�K��֐L���}}��U�U���N^	��n����Gyg������aj|T�E���L�^F6����w��x|��U��K��&�9F4e�ugd�O����Y1o'P�1���zv�U������3L@���EU���ԡ�� ���#v`U����w>bO��%����d��t�u����������t@qFM\�U��z�'�ɓPkS$Ov��.�7DM)�w��8�&U7�Ѐ�w`��_�	�W�$�)C~ә���L �������[��Kc�6O�&�u�f>�u
z��֋a��nB܁�խdC�DY>��<�d��q����|�Φ����L^2��3�<L�~�{����!q!�V��j�x�o�2�����t����$�l����g.a0�����tr����4S��ͫ��!�u��6�� :��YE���q�C��YF�ġ̣�8�)��T�7Ԇ1�5&`v��܏M��17�����}����C���;}G02�B��M�Pv6�"���� j��,Ў{�hq��%O_��Qރ��'��CDDZ�'�7H��~?��y4���02�R^���z����&���Xߒ���M�$�7w��V%
��c]�%��?CV�ړ�K0E'���,�y%U�K?Ԓ��#����T�Z+y����-���H�e��@�	�����5�tx Y���N�[�Uf}pF���b��w����e�(CB���5���DL�9�Xė����mž��^K.B��]���v��l<���x ��Ý�>�p��폯�Jc����$8����>vA}��X}wN����g��w�O�q�&�k.L�@?�ll�Eۈ�zR�'�y9׽�1�#3�~�p9�^��j����6�e|��Y��N����$���_s�$�n�x���}t@W-�[�w�9�b>��"� H�LC�if��^�j
�"e��-����SA�Dԡ؜�D��� �`Ԗ[�����Schq��%-^�k�M�����(���t�&�]u�d� ����&=�����ŰΖ<�,�pD���T���9�O<s�I�+�,�a�|(6���
R��P��Nc��lŒӟ�����6�D`.;�ZJ��(!���Z��Ɓdi< ����
����L�Qp�������β.w�~�i��4�/��9j��l1ݞi9��ēԯI�<W��t���NF��?�|�F�@'����pL�pqڙ�bt�k�Ʒ��
��~�+~�$Qقu�F��lV K4M+,�b%�n��+��ֲ_jjz������{��~���ݳ�׍�׵Z�|����94\�X�Eä����a/]�{�x�ulD�q��(�T��}�Ἒ���BQQ݊'Oc��R�
��z�����?k��ρ�����6�W>=�����������CJ��R��7����w�"~�0���Ҥ�=��Q����Fě���~s��N7�s>(;�1���258��Q���K�i���e�hL��Np
�Bᆋ��
�Y���`E]���p�/�"�F���! �((���%-a᭯�APE�vItH+mw^K!q.�$��d��d��!+^5�]�m�vi��AC�] '��nw	F'浅��t�v�ԅ�ƛyh�&e1\ԯT~k��S�&�жD�DTӴ\�⯷y�o&�V2��d��������5^ M�V���jM�x��/��������B����@���'��7(���\q8\M��������!�C�Q#�����C��ڰNo��]�ߘ>R����~ f7������E��5Fm#"�R������/��ڄ��Y^F&À�m�_;G)�oS.Ấ=��0��,�\���t�����F���,�WWE���Lxɸ�u��B� 2U�'Y�ՠ�������/h��5�[W|�Wr�xN.�Ic�Lp:��/�w��Clv#y �tǈ�֚Dč�U�J�U6�$���4��D��@Բw����ھr�j(�8+ ���&��K�5)��k����j#4�4h��L��g�5�DPQa��Tm�����bľ�9&{~~b�&�c3?To��&z�F�{sT�I�`l�N�����g��e�sR�܂�u��p�HVa^֫���bQwU�I�Zxw�3��ֈ�؅�7\xn���s?��
�5���a�u�~3k.�l�tZ]~�z&�TY��!�a�V�S� ����cV_�l�V�[o�ׄ�|�1�u��5T��qy�]���8Z5��|?�
�@/��6��S69���!܎]b�M�pB��:AP�*c!�`��4��4���;R�n԰�o%��1�T�����iY��~��.)������ �<�\`C!:��������+k�%M����͡Zf�x-��-WTQ]y������յG1h�p��ΧS�y�dd���wR�+�H��6��{�#��'��AMb}�p����b�Έh3�l$!#	���5���HAY�O��B.���(���f�a�{0����?��ƥMϛ�x���ίO(r:J]��O��7&�Ida���'�M��U���5��{���Y������J ~�)�����s�R�^�}`�����8y0s���6nP���L����o������\��)�3Pk��� fa�"��؏�N�^��̔����|hSt�B�+;U�\��X@Bu�*yϖ	�	�;	�f��c*��ak|,�\�?l$�����H9�g�@�%{�ᯡsА�3�X5�D��~���,K{�u.&q�v'TUn�J!����Jbε檕(�L������@W�
i2+m?��� Gʏ_xҔ�K�C�O0���P�`'.��i�o��Z�S��ؕ��_j9�
/_��Q^���f�bWI�Dd���.�����KK3��T���.�4���L�L�K.��@�L�����"G�����Ә��m$H�O��z�BsD�c��省)V��7{5:�B� �7�]Qf�8J2�3+�o���Q!`�UZ��U��)�f0��Tݳ3n�+�+�L�l�d/h��a`U-��
��s�L��8���L��t�#O��zB��Qv��5Q7&��������L�`
��㱠�0���A��`��>��٭�@�0T������9$�5w> �T	N�+�vi0[�0	�C�pZ 0����Ny�j�;�u�uf�jguh��͠J�39�2�CF��zb��!�Fq�w�<X_yb0���0InB�4��S@��J�8d}�D��b�4v-k�O�P�U`k���s��lqO�X�L����Q�֟��0@��p���9�D=�CB>��?Dm���֜4� �8��YgL�]^�ys: �7T!g������4��W
݈���*ER�bIE�V�:\��M1�0�B��ѩ��TjhO	]�B�����noS�ց����91�nɂ4�`KRFp$�nStU틉yt[���lX�o��nݫ[/8GFY0���������@r��2��"�#2o������'u���V�]=]Ehb���@w5�m)GВ�K.��.��{.�����f�%��)��_�S�S��$�}%�ejUHw����uPd,V=�-4���2�28��X�כ�~��Λl�&�G͊^��iZPj�C3��	��;?�j�?��z��j�x��B�Qf`�	rvI8�j�;W��na�ކ��#E��ٴ�Wԋ�d�P���^{�^�r�o��k�|y�f�'4g[�q�;<�Jw+�����!�W�����Ў"��8Q;�ڃ�^�W�ժ�4
��B�Eoo�A݇�b+{�7?v�8�f�;3U^�+( /*�'�n�5Q��*t���^� rl*�D㨿���K֠�ؗs�q�z�4�T�d�Mz������K�`�^�mlEu(IS��D-�F���h� ��IŢ�cL���鉘Ӛ���?~��=V����E9%B�ߑ՟�+tb����(�ڹ|�6K9�dj!��l���*N�@���E��fPNu�#PJf���t���]6�/�H\<�I��`�q�=���.Ys���h,��0�,��i��V�Q��WUn�� �تuB7!��̩*n_R^7~v�3C
F�=q�	��i�+�h�q��	���TZ�ziTN� , ����e��FX��I0&Ch�Iά�R�^b)|����e�������<�q�x��8���s��^�w���O�1�u�Ц�^��X>���W���Mw�B>�.%�^�U�77�iJI�Ӷ�U�R�N@9�z��Fj�[[+�l�Y�eo�0�V�Ad�b�!�b����ɍ�z�Ϊݹd�"�s��U���(�-��y���""h*zE_h��w��Q<�8�i�x/����똜���Im[�8��ek,̔1�^�~+�(M�U�����K?�J!2�d�>�Vi�ۙ��Œ�{��O���P��Y���a���'�9<�_�Mv�N�r���T���(l�Y9��J\�2g�%��?�E���leL��غ�/7�|b@tz����Β�ǆ@�.
����K��wFT\=N/-�]����]]�{��@�&�Cn�V^u�8��US��G9_�Ok6����O�x�`��]X��x�fB�vᩣZ'4v��\ӊ�̏���3�͈�I�*��NF=0��rrM���4�\��Hi<	�&
i{2sq8�O����%L��+���#x�HdPM��"A|��:�1�d_9�^z���& &�A�ZO+��>C��HI�C�i�fd��ZR�Mq�j�����IDP��ILȮ���rI�_�ޮ����1��z��)�T_	t��П���v)���YA\߷ 5{�S5� �=4��?/x<��~�wɀf12��q�G ~�Ȇ��]��̖̱�nj�"nr��*}N�x�n�6���1Y�.S"M�;�oH�B!�J��K�Uy�!�ye�R�b~�ly��	�����T�t�;C�"��*�\oc� %�bl����rQ5q��UZ��Z����N��UΈyM\��V�7u�v�3���a�.�1�_U�E��d�Uw(�ӂ��kw	/�\�;`��mm���Ą�q���k9;������a>�7�Gp�x��_�q����J�<���ě>���$c���|pӜ���8h�I��+j��%��]�F�J|X���x8�m��{<�70d���.&��3������22h����OZ"e�8u���/"���	�4�y<�_\�n1s<�ߚՌ����ө���L�t=y�֭���������J9 �aF�Hy[^}un�����WT�Z�k{������R�TϾ��+&����v	�V�Ul"1�w���tmgTG@���CU���{���9pß�o�	dG��c����颜	N���u��Z5��0!:sp���m/��C���kQ�JD~ ��C�'�5�?-G�
H�g�ӝ\�y��6�myI�1�*��n8���H�$L�Jo�o)�# *$���l/9�W����?c����yAv_��J�mt�8B��^x����߰��f�{��_N{�c�)q�D`���K���IiYgצ�����E�������]İ��CY����:����oP�Ju��(s�D]t�5�@=�ʫaC���%�@Y8�~}��@/������07_��л�ǬSb"���!����!zk����g^��B�ᎉ��n��i��d��џ6�h�˗4����$-���	s	�_��L�	��dD4�
����ď����Az����,Q�cxu�yx|�W-�GxI�X��}�17��)��铼�$`V%��~e�m���1R�"��Ԙխҝ/�����qc���_H6�7��s����\Ǳ�W��,l9G��ݳ9^z�n�ͺ��@ꜿ�*�V�B�Mj{�'�ZZF�q�c�3jp�[6&���W6kHқ5Zori�[�a��b�"~.�Kh���<��m�W�=��Y�~��$�/Ǽg�pk�~o0����M[[5��?Kx�Y�h8�?���8Qs6��߼�+���%�����rqf�V�j�wj��/��X�Nieu��D3���?�d$�	��z��G��w�37�w3��T:,���˦a��NĀ�[+���eN ʺ�D��=}5�@���[yS'���Yv�Pԉ*�����N$�LJ�~ޖ��Z��{�X"^��������/I��q�~��V�����g��^��td�kED+��B�|�I�M�V�و���w��ݒ]g͗%6��C|!�z�p������x���,�C21q����v��pz�o���Q�ppR�W�Q9a*����<Ӆ�z���lp��f�ABX�C���·�IW��`�8������	��+����r��)���h��3��q4���Gj��a��$��p��"�g�/a�[����� 'a^X�43�����!��Ro�\���^��B��;�0rü]r련���lTp�/0�������A �\ټ*M�j*q�I*��U��	��Gpax�aK{�j�,�� �xב�c�u��Fe-�S\��BS�Qr`�ӄ���{ՕV��x�V�t�}�G������g��tG�@�N�^� ���3 ���	m'ç�H#�Խz��G	�c�h��oJ,���n��jt��YdJyvL R�Y���&��G��%���B�+�5j��6����	�V�,q�њh#�@/���ֱƗ��/?�,\�u^:��"�������5Έ����غ���έ�}�����|V�*�UK��m��<f�C��y�u`����GIjp@o ��6�M
�(��(�����7La�Mx���ur�*e*R��$�p��İ��++�$X�Q�fk A�)�r���B���Guӥ�fm��YA�@�#\;�>���K�I�T(E��zr�Bc�cUq�T@7��<ǎwM�C{��_��0;s`&�֥�}���5b���0k�(��#�g� 5���ct��Cc�`�&u\1fLTY�٭{��x#\C���|˻��o���O��+��rs�{���HF���X��u]��Y�>�珖�;h��d����BOU���oJ;he�?[�w:$Kb��A1r�oa�����TH�l���m	:��dx�siqH��RV�4ܖ�ag)i��6�.t�ApPݥ�ޕ&"ت9x�R�"���k�hr���̙��;�r�҈Bm�Oɲh�
LY12O���[̠S2��e�b�&��ַ� �����W���Ҹ&l�.e?�k��{�Mj�m;�ND�xh�-ҁ<z�e��Dh�/�ħ���HV�%<�0g�2ƴQf�(s�y���X2��.�e��!ų.�`Ql��� ����
̋���tS����cG�G��Q���5����D���ӛ�*ʀ�ic�7��^�+�����	�=X|�
��jI�RՒ��B:��EW({�gk��KͷZ|K��L*�5Fm�F�}f��7{$I4�P��Ϳ������$��W��.��'���(;Q�d�^�@�o9����|�v��d�����/~0ؿQp|�	����!	��`I�m�EK!b�C��(��_�?r@���+�,��:�(W(����H%��ygZ�n�X=�%Uwb܋�f�v/���t��>�z,�DE��oh9s|�%,{T{���K�����f����Q�9����l���{"y��>�(�I��@�jA�q�'��D�/�٪:iX�S �A�힝loG!��f����0-L�;+��E.��Ը��8��<�&��67Ͱ��>q��'s��\�h,l#�d����Lj�Ss8:����7�+P�J�υ��>s�O6�B��!;�3ՅK�(�������ȌN�0�&Q"L"����N[�z�]Q��{Ń;�����zټ7����@�W䞫�u-�E0u� ��?>C��k�q.�h��# ZWkl܅� nǆX"��\֌�
S{|��F��&���Dd`�Ǌ��1��&Pr\��F�<��F�g�n]�y��cvԳ`�DB���3&�ʄo�8��p�sJ�Wĉ�\\�(%���S=��HZzZ����0q�V3�M4��w}I����e���}5i��Y~�>�}W��
�:�ո����̒b4J�b�E(}���CB�����;{� e@���8S��f�Y���{����BpD[�D"�qjlz�C<2��w��Ȗ�����`�}>�R���n�:O�:�ǡ[X������~.�)K��Q���*��ތ�q�9��7���pU�� ��6��t��4qss��O9��6r2��ڌV�=�ш��e{(�H�G�I�o����~�>��8Zc�гך �X� ��
	Xr���[u��ӟ%-Q%j'��J� G��P�b5�[W�!��#Aw���������
-o�R�z�P���R�[�#H�W}_���ŭֽ�V��kr=�f!��~�gZ:ٹ�UͶ�A����ۀ+.}�]T�(.�U���z�H�4΁�;8�K�6XR��Z�C�5Z~5"���+�����v
p&���s&g'R��L�	������^!W���÷E.L,�q�w%5����-��sK��E�M�~�-�! �g=$vC�D��4�L;�k��f�oi�c��8G��4"��WW~H�ZEH	e]h��e�a��<�s�S��������3#�ͨ"F��l�*���q�&8o��> ���սW��Gs0ȸ�8��P�m����A亡�����?���?��_T��ZK�`<6�"�)��K��D��P*��d�NZ9���@��ݮ�3����'J�<v��AO�Z�"�$�(C�-c@�o@��H������n!��� je�M��jj��ڧ.	�.|���R�Vh�E"�Ւ3���_AYC�k��:��I9$�ԶAT���,�- 8
d��+G�ƪ������(�����PU
_�(�^����0Q8��{�XO�:���v�`��h����d�hx�92$:w�A
<]��.Jm�ꜻ�����������g�L��(;7l����j5S���cy_���;zY,7Q���甕���f��/��'Ű���&H�!�>a���ǅ�*��܀��P���\"cb���uB��5�] B�c!%� Y`�`�To
�'�g'H3�����,��ו���~JШ��[O�e��^ʏ�u�8幦�l��Xi~5��O���v�k۶�n5����D<��<�Bg���}av��5���y��]L�A�9:�s�ㄝ�'�>q>m#G��C&�P�-o��8�1�z$42��~�������T�k�	1hx���>%t�_�h2�cD�u�}#���Ŀ堏��}����B4%VVX�|�a�y١����G��L�߶jn�G�`J�l�<�
yl�M'3s�RG�K�̘��oݧ�F�D0v��?���*�Ӵ��â �7A��VKn<K�hC3#^���aq�Um��V|�E��]��1y����B�e̔>0�+�g[�@VL�\s5"v!L�>�K{yO

ed���%y��_u�1�PSdϽ�0f�.���J-,�a�r^�ۋ �s&���X�E�@�;�r���G����!�Ѐ9u��\\��+=�����ӽ<�h%�?�����1YzߣF���\/��^�����k�>x�q�>!�A�Yw�֟P̷�A
u�^��e�E���o���Lc��Y�M��稥\q�f{�Ot��	��l1 �i��t��W�р��W��47���|�͠W��z# �ӵldZ6=��=�����'��D6Hlی�"���|ڵ�ӈh�H���ϑ�����l=���dah�\�b+�Ƿ�����h�B�&���6I��2����嵍���N�z������/3G��J�ց�懨�-�L�.X����f�:��si#,�vr$P�&�S��6� ��bY��� 
U�Z�çݺL�������fL���z�sӫ�F^�$��X��5A��
���w���H����{���TH0X�]����<�Í$��>�HS+��|�rWR[	d
"��"#���͠��Cd��E���#X	pj�#���K���m���Ot�FF���(��t�"��(YZ�s�m���w�ԓk���R��H$�&�#����7{3�Yq��d� ��B���g�M�ˌ�%�*�mv��qh��ܾ�����d����'/]0Q���"h����^��ё�qY�a9?���e�t!�Y� vs��5m_.��W��!��y��/������)�I
G)��Hι�N�3�ъ�
/�f��\8�3ױ��i��#�F��c�}Z̐vr��H��:�A���֧
Dz�eu���+OC���ל���%��8���}����e��o����<.�ܙ)��S r頼�t�&a+���\��!���nQ	&o\mDd���I�ИK�F�!������8u|���0�5R���]ct�A).D��e/@�b6K��?�N�HR_���|v�C�}�2�s�M���E��Qo���,����Z+ܠ�k�;�}�����}_�Κ�;>��j�ٜ����e?0Nh󦟨�郵"��z�&9��u0�o��/�5���Q^���s�80�;0��x��M\~n}��p�����!��=C��Ѯ��R��3�N�!$)7�zC�L�J{�~������!bg#�,�^)�#)���^k,�uV�Dj������b;W�.ߺf��Z�bw�U���&X�4;��O^aV��8���t����@�̷q�~�L e�Q,�k���|�ܠ*=���/~yR�*����u��U���4�@�w���Ru*V���徃��|�i/Z/zh
������x��	I��{�"mY�s��	��
VA�ݼ���	��OQV�f�ū���'�泚]Sx��n�Q05�K��|��&�w�V!ڷx٨���5��4�+�2F�����n�����]\�8����-@I�hcI��3��^�^�"FjgR$-��Cc0��_\��)m�.�� Jq�Ύ�d�ul��L�f���Z�����Di����6�n*�
l�%uB�;�(�݄�ގ��{Ƴ��+-����S����[�"�cI
����"�[��?��)���[�$�y�s��ri��K�Gָ䕅	�UH|�K^1&O�#�6�!<.��&p���4fû9hZ���<T����p�E�@`�Tw��"�m�^�>X��\&QND��{�=r�A6W��~^N��7n�k����i�7M��g� J�W^o�r�v�, X�
H D�31CX�^&x�M��g�a�(�;;�J@�f����q�r�ri� {"npQֳQ�Ih5�"�NDdc�.'�c�� 8�
̗�Z�i�{��z|#J�
�	�8���Fa�Y.��+�xb��	>M\o�\��3�T� ϥkL�a1��u�H��щ�M�!qjM6%��s�{JR=S�\����#s�ȳ$�D~���i��)����E��`�ij�'$3?Z���V[N��6BB+����H�\]�vgƏ�EG���D��� tY��_�_|�>��>̖�a34zҍv���x<�.{�4N�&�sCUՅ
m�tG��c�XE�3}U������?�CV���d�]X�*i���
�g2��'s޷���P�1�6�*MI��a��oM�"绌vC��
΂�శ4�ϻ�� nd��`��
C��2�q�����:Y��j�[E>1.���	c�Ώ07�1��h����l���  ��Aa��,�z�;a�Ao+I��/T�������Ox��N��e��:�/�CM�I���~�9�	8�p&ʖ����_E�>����t,/�Ζ[�&�0O/��7zV�i���K`/�)P/��4}0��RmϘwc�)��p�K�yG���(���:�WɃ���|L+�Dc|�Ej:͟��N���U�#����H5ߞ~�	�{��8og���ŰC��Q��?����Z;ny[�J����_�ZB�#��J����"��D���{/�o�CT������&/㾌�h�,m��"���O��.�@�����Ng����C��)]y�T��
�)�=^�`}��	�H6r��K<u��q�G��9�0�{# 3SG�.��}0�f��"kY��!�}'w���E��Y}jᾈ:�8�J,���DE�������ܘ�DC �b(6ܳ<t
B{����yOM��T��Ko�����e�� ��Ԓ��T��J����?�I�(�Ne�$�߮����GY7���1R��>&^Oe*�s�j.w�'5E�K*���I�g��A��
^lg�U��F�u�A�x�č�J���@�'��� ?�,���{Ի�m_��#��rl����gf�-f�<����hJ�'�͒M]]�UF��1�j��pG_r���vP���B�H��h�Ӛc�u�_�}X�����+��R.�n�N|�Ҋ8ta���0xE��[���=e�����̓��u�]��ta-��^������(���j�ۺ$�g��av�u��Uخ
j�^��C0���I�x��d�K�t����tRNA2i�4f�ܾ<j����5��2 `)P7E(��q���iL��p�@�r-ӓ[ �F��j�!�=A

�MiO8�$�ϓ硰�Npr��+$8���̇������a�`o�M5(�r��Cт�ә�Yf�꟔�Q��6�A����ȧ�x�r��I�-�C�Ik���a���ECLG�W�#`[�';}-�x=�z �w�n�P���lT&�t���4/ E=�2�=է�ʋ��}%�֎�d&���bͷ��"\�s��u��S�90T3�M�U$K�V�[L�q۵��F���
���y9���Г�׮i��݉�μ���=��uM-H0x8�-��������q�B�Օ!ϱwe:	��*���(a��+L/��|�����i�Ȳ���=��b�q��PXQ�`SV0�[u�	�f#*n�V@!��W�q��pK_!��09���e`��_n�{�����GFw܅Uv���?3. -l����;փ
#���x�?�3H�6���%����X J`�Q��_��W8a|�m������U�TI�*�&ck���^8U ������EC�ʠ��Wd�G��X1ZjȻ[<���!x����#{���w���3�'S�"Z�����>��(6�4��#����\?�J砠f�#������e�F��`����0�a���,;�n�d�
����z�\��@�������p����}:\J1����xBE��z�J�|�@B~�X��C��$�%�>�z�p���'�HQl�0T��J��w�OR�IE���s��%�]�3T���|� �2�H�f��֎U�VB^r�����zc��W��9��ը���x�����S�
%N#�{9+k#�YM��գ�
���X6�e��q]�f�����(כPS|�������i��!`�^߱h��|��r�!3e)_�RW�&�3�,y�=U�Ä��Bڍ;V}��'g?]��ŏ%[��]{o�ͧ=�>��{��3�EgEa�D<L+�/LNXd2C�￑�R[�gb=��MD�2�u�����C;�j�[���C��C�np�ߔX�E���9��=�݉����^����8<HVC�jS��J�l"�>*:21�0��H������۬d��)n_��uj.�5�.�oB���3�,ੇа��K�ە�����v���s�ɜ|u*5�t$��+����}B߻?��&[�?�V��+�)y!l*.�XL �M�92H�4��fJ�V�e��e����#�Ɖ�p�uM����{rh�N:���Ԝx�`�Q�I"�8�:r�W����*ڌ]޻��K_��ٍ�����Bn�i�#����i��GA���v�G��_Ǩ�����'��W�#If:A$�h"w]`wO��u�ܑ?�w!�j&kf�b5�C�^m���1n��چ�p�ؓ<f0�o�$�G��*�XD]��mR��΢קk���FŶ�9����/ES�jyV�sE���6���_���VQh�]w-f��?W&[���ΤQz
�тȒa��K��JC�g���/Ҭ= >�K4.f�o��G�� ��|P�z��Ƴ� �Ҭ� �IL&g7�љi�?c��E��KBi�����m�v%(�*�E�K��K�o��������"d��«B�7���x��|�&C��4.����w�5:���2�ý�O�n���ci?.�j���G�Kf�ƥx�uy���hO{���h%)v
�v��D�5�?]��MnZ ��O(j��р>�Ź;��^`o,B�Y[�I�
A�c�p�l�w���1ǂ 3�PIp�SR	V� �)<+�4�{%����3qOa���H��>M�2Y$�A��K�.��w��rۑ(��pEqK�0����Q{	H��q�˝��3��o@���n�W~+�s�*R�e�!~����"��B N?d�}�8�'�*Kh�>��:[�A�p!ri�tXT��	��*�a�=�j0o����.WA�O��/��ŭn�H���6�7�ɰ�b��9PkWIFѸ�[ծ$Ǹ��,-:#{�<��lI�ZR�ա���y^��YG/�?� J=��	�8�DJ��`[�M}yJ�Ul �z�#uq��Ҷ	'R��d��,�s_qʒ�o�E�`�&^���rT��k�� �&D��ʊ)a��g�\[�m���MTV}7>�F��Q_(�?���Է�<R[2$5&@P�B�asV�O/�`�< �0E������eok@�;S�%זN�6�3э��ɗ)�b�,��N�g��c��4��%�''|�֊����돬	p�'A�7�ǯ{5ȥɧ��t�E�Os�b��g��<���̸�%��~�N�ԏ�\5-Q~��*�y���.�����c���BU��$-bɉԒ�6.���9�A
��/E=�q��_�G�͸�[K���L�9�t���&)��v�P_���Q݃Ye�4S#�n	dMudD�m�b"�՘HX �,���r~Pи����������l�H����ߚ�;.����:���Igw��ܲR��ң�X$��L�H�|���w����<t�R��d'�����$�L.�13�y�?od�Fr)���\u������et E��r�w8$���a0�D"�W	�w��B}��G- �l��4��o���1/҃�9nu��������#�ݾ�@��Q��֎�_�P�j@nǺ��!�K�W.���L�B�>m�#�|X��l�;���R0�,��fFD�
|k�؆��HV�'w�byd�޴-U���'xa�q���e�>�a��>�ɪP�D
E�SA-�O�x�����Sx��1nN(�6��βe	���3ݧ�~H<�P{�=>��ִ��/�h�G�[z�e>��MH����Ɲ&��NÑ�\�,��J�ǉ~���݅�)��a�l�AZ�[NQ�~�c�Kh��q]iF��<^r�X�N�%߁t��1�vXj����gxn�E�����Y�-a?�\�^�3A?���\��Zdg\D2��[Sx��z��!��X���l~��O��7W[�Jd�]���sG�x6��'T����C�y@"6����u��k ��ݎ���/��Զ��e�d���݅�=t��ֆ@}��lN���zn���%g��R��qQZ)�^� ��P���LO���+I�������b˭)�h�H��W,�h=���5ք���)�h��ť�0�(�	��0��j�����7�� !+]��[T��ge���zWj" ��[
ն���c��G�&�����2l;�H�t��~F�=���ަ��k_�jp�=�y�I`_nԔ"��*ǖ�z��;u|��(&WS&��Kن��Q�Zy��:=�c]�)�*)�����K'MXKG��#N9���U��*v��v�d.;����H�&A��8ޗCg��Í}��>V�bz����G�0�>��g5x� نz�@�錝X��w~b�7>�܅��ț����z���0��[�Mrq.έ���u:�I<���-� $
���#>�ߍ�ܸ^c&FFF����7�0IG���yR]R*��*�e���%�.H�N�<z2�F����|h�>�<��}�A�Iy�^�Gcʇl�V�V7yC��h�U�IC������ν��z�����(u�)��6�lv����
u(l��ڪ�b��B<vi ���W���3}zU�m������ߍ�Y��"�\r��@y5S9�i��⾉ ��5x���=�����L��KH��ܾM�^���Q��]rBiG��� �E<���L#�`�zr����U�\��0s�F���sM=��Q�e�����_��E4=ޚ�A��V�M�l:�����{N͡�v&uJ���k|���5�k���Q���+����Q�c��HkD>��Z3��,o�񆕥��L^�z��vv�؎�����] ����D�~F��A�3PX,��[�m���bC��,�2�����{j�_�a;)FRk��?s�lp۪RƐ��Ȼ���z/�Վ�p�`��,hUP1<�Z�¾D�ќ
�M������4:�cq�=}k�|�UNl ��{�%�z:y}0"b���y*�T�zaa�����tʌ�9X�4��x����[�s�d�x�0AGŵ�j
@�L��BP�4Y�O�C1G弭�t��L�kB��j���e0��+8��i���
��KA#O_m�a��y�j|���c�%�0�+�	Q�.���=7HlL�M���D*v�m��c����
�J��]�)�w�=����+�a��`��\7�҃*���&�c����P���2��T���<? ���V�Ћ��ASٮL�1��۪��`��cr�����ۧ�M�וU�"� �+��d��>�-01���D�︾%�JI}����]�Y\��Ssq��I�Ǖ�I��`Ώ���� �)����g��'��3FG�q�G#�K�yH�B,[<��H���/g����
��ϴ��9E���_���N�F�z��\�:TX��[$�=;���4��"�r��"+(4�ͮ�Q�o".�������8���L�t��<��v����k��j>�%z%s/X�D��ºc�[HMàl�z_&�>A��Eh��XV�JNrw5�p��$�|��.!HC	3ie�����:�z<��3�/Ԉ�+�K&FД0-�%h�B����",ܢ&��y�L�$�qkii
pg����.�e����]CG�眇�QM1T�o�\L����c�i��*T�z����z2����U�q7'֩+�;��͏ ����si�.��$��S	}���dޖ-�s�ùz�5�T�Ȗ��j�����.�	_&K�e�����`� Ѵ���6������d��9WZ���d�6f���+�΂���Ɉ�ҶY��eh�}� *W���#�>n�����c#���|7
��]Y���Ɩ�&)KA4�>�W3fL\J�Y�j��`��5,�b�	�����F3!ŵR���7����Ո~�[�ƛ� }9��� ��Bd�5��9]�Ԅ*� �I��!���n�L�o�p����&�X�:������Czޢ��݌�^e��(�z��YaS�t�WL�B���Pސ?đ� �U�y�]��h��C]��qW��u�٦��둾U�7o��h�T�����0���@�����''����P���V`����U� �����Y)�㌓!�~���'b�<>:o�����`Y;`\t�z/o6��As��,�<N:Yr��Mo^&�yN����GG�_�ˬ�Ӟ�+$�0@�o�,Zy �<.�]��PGg��m�ݤ�FH	'#���=Y!��d��N��4|c�($S��Ew��u���2e]�z��r��N<�olk��g��fr���&�&a�8&-B����{�|�:�7���2�t����>K���]1ra�xn��S��P��z�M,�k��sXKQ}���@Qp������S��)'O�v��WξK��Z�Z� ��xc�������"}����~t;����S
a���|�0^e�U!"�08�L�2���s%t*
�&A.FO���_�C�Y.*����In�!��$�4��%ʽ�=9�}�?�߀��l�n�WX�?�7c������6XNFJ)��]ϻ�V�[��1�� ����[�4�ᗺ1قp�X'�'6��/��'�2�Fo��(>�v`$!��)�P�#t�2Hx��h[[��B8�'_��ұȾ�ħ7F0d[��\�|t���bÉx�,�_Z���5����Q2����u\@�Vⶒ�6E�H�@a|`�G�fD+~�m��]�!}�ɹ�f���&���%��D=�t~H'���[0J
<w��L1=�t��_���qCX��>Y�g�u�H|�^E���|�������$2��X+R����褠����A��L2��y�h��`�[��-�#��	S@V�nrb���^ ���F@��l4΢�Z���H�\a��>q�ǻd�q���"O���������q��.yM@���d2�J�%�\���&�T4�P������4z�]}u�L��z�i�N���׿�W%j�G@n#b��|E}�P�`��W{!L�!�my3�?$n��Am<3͗Hi�r����r�~2lW��[Z�PfXjl�O��׆f(	U������ZӜ);��բ�ogS�b�pvb�a�ԛ/Z�OcY����'�5�A��{����%�-�>�x�4l�V}҃\���p��`@U�x��&e�N��^�#\0q�W�9�%?T�Lk�]�����Q��'�OKD���s�!�I���`%�г�<�/����㸦n�1�,,s��P~�:՚�.h�GIE��\����p�B��c7b�~ZR���0y�4�p�q��ch�� �[��n�ԪN�x�S�7�(��;O�u�T�"��P���d�@�@O׸)�D�lB�}��oAEh�Z�n`�2L�1�Ǯl���ݺ��O�����gӲ�(<6����p�b�O龩 1e����ƨp��-7H��d�j�����k��m��u�b k��B/�(Q>3(�9_/p�u3�ò�J���ó@V��Z�K��������&��&��ЅuU�#)���F����?�5�e��U�G�քu����NZ���PV6�)��?�h����@� �R��I����b鞽a�������1��G��m�I�'������<*ӌ�Q����-�i�u��q7s���_����hg��f,zW8
JyM�Iv�8uj���R"p�~�,��۞p��̟�a�Ŀ�y�ub���ف$0� 2 Q�ƴQ�l�Q>rP.�/��������"3� lXV��&�q��Ջd�"�*�0b���o|�B��´�DS��yR��&8�7B���t�j93YB[( �ۀ�S�?��G�B�s�� ���,:(�&�U�ļ�*/8<���n���=�d��I�AiˢIF�7&�9�jP�ԍ��S�ٴ��^}>�0���0���e�O�qeP:�� �*��7��݉H�7��p:��.X��XV+�ڟԔ{�l��0l���b��"#�l*ܷq��ȟ�����v|�/��9�������n��C�N��͚�����с^0X�խ#��DM�;�NpM!:���B1�1%1�*#5����d�f��Y�S�d�f ��_��8n3�
"���rIY�?Ƥ�2v;�y�� �H��FY������-���)YT>��M<	��PLD�*��1f��ғ p�N�!����Ϩ���#R����u^:�6A�\\��eo���:�X���r�|P��$���k��(G�%�sr5��>_��N���^�QDIN�>)��y�c������(�O��d���]�e����~�]��(�ϴ��)��W��H:LE��Ζ_�Ga��ɍ�zփ-�S}�TUNI�
�X-V�;���V9pf����e1���Tlj 2�5���*:݁um��ϭ.�
�lME4��x�|A��n���{4���n����Ȁ�H�O�qa��Ե�V����|����
��!��m$e�} �5u��ƽ�F�����`ʭ�(f�<�b�~o��[������旾��5�=^�N��B��U5�w?�2z���o*-"�qT���M�j:�OO�8�9)��uؒ�E�}�` }%1�0��UнY����볨R���D!��9�����c�?0D��=x}�V,	P/4k��S��xv2�n3��W�w�B�aU,���/>OxA�ǫ�|�g./�UJ3��M��dQ��P��$�˨���� ��@������Y�gQ�z��{{$26����$�5[�m+j���_ ] �P:���Jΰ�xiRX*.�PU9��]%KLz��W3��"�h�dbI�!(���K�uT�?R�ʯ�_
��P�`(��+��%�ek\(R,\��HZ���i����5<	���պ����9��n��h�����;ǩ��ke-�"pSx���M�D�O>ă8h�7_�*)ũd�<��p���g
6%��\f�!�ƵA��lK��
V���FQǦ��+�5����q���8�a�)�*Ց�b��U}a��j#��T����N���_F^m���󃯒7+�&��w^�������F�b}��'�]��g����������dH|8���K�`�<�5���~��)k{KS6 3�'�<D�V��ը�>��Ҫ�ny�K����ۜ�Y#>ɯZ൓Dj�/��Ǥ����[.����GoH	���>@�L{���kʩvk�z����@�\el�����.��K��jw��@[�m~1�%�$^6Wv��Ò"��Wu�k!s�gŽ�F~>=~�*(�.��ӻ3:�j+v�n�8�r�3]��t��"8�%�v��ݐL1��`0X�K�����o�S�,{��X�r�����nU���[�<��׃��Q|�K�0q՜�����9��.�+�~�~�����~X�F���ϩ�O(|�3�?�+^���\�}�FAʭ���֠�R�C����i��^�e�(# \�u��2�b�8.hp�j7�t���`�z���:[#���J�IÏMt���1��A�g���2�{%�-rx��fq��!Oꀎ��̝@�2���Y`	�>�
\]�@��)_�ۭa[�N%�٠�W��\|�6ߧ��]�]�um����Jo�����Ӊ%�"foxA#��B3��R��>a��?I���C��0�/ٮ&��t��oz܅��A�q��p��3Ǣ����eU��GU5q�meW��bS�P���o~�l�n/Z�/KV�^�㊠o�c,֘�;V�(�8$_��{%��`Z�)XrImL�7.1V�G����Is�N�}8J^ፘI���\Ǌ�6�F��d�F (���w���J���#�:���@"�ȥ0��-'~x^�	�q�FFb+�Fx���@C�uf)�@�֫��A)�>+��'"��5��� 7$-�,����(�^+�$�i�ꃳ�E/�	c��
�v͗i8@��3� Q�����h��h��!��?�x̞����`X�-P~���U����f~�x��p�;#�}J�%�<���������"�G�&��J)c��<�@A6�p�����Fۖ:�8�9��(�ޝޣd��Jf��|���9�����;9�p��O�Z�	��5['oN�)���Tf��o�pDV#�6U&�d����迱JG[G/��Մ��OɃ�hp�'y�r1!����/x������� Z_ؒ�� ��%����=S��O����|�	Ed��� T6�I�"�J2k��mDp�A,a  k=���+Ѳ�4l(Q
��m�Ӧ���%���h|�U�?�Q���fݍ�40IL�>�u�W.��TZ%��Nj!���F�LƑgŚ��պ�=�8C�
U����j�Z��m���~g/�Ipb��� �����Q�h�9K߮�/> "A���D!�Y<��)x-tV�Fkz���Y��f�K��g@1�4L@J�1�Ǚ��~�׈LA����f�&�Tp�;�z6`�t?��6�X����SQIOm����f�����@zV��׮4����'�^Sv�3�����t%N��#��7u�[zC6h��tee�E$��6�N�ETN����ᜌT\���C��e�}���.l�٢��;����u^;X�6�h�靌/��]A���OZq�N�>��爻)�=Bà�zKa��l���,[p��cp�}��Ӓ^����vB�R�y�Mq^|a�!�逆��s�P�N�����_�򕜙x�i��� ���^AC:�IGOϟ�"���i�z�[\�$�Mϧ!:-׳V�}�D������Խ����Ɵ`��Y�h� �(�R�	�ՌX�'�W jO}���l�C�<n�ŏ̈2 l���� qp��Cm�H�r'L�ZP�L����5�l��d������XY��&0�>ጼp5���;�7>՘�e�ڣ��4����	O����3�CRV�D&9ui��k��,�S$K��� �[R���߲�
y24>�:�����i^~�]�o���;|��
^��Ώϲ�Y���I�Q{x@O ���|��Br��r�[��.%~��($�u�/�ҩR����¹�Y̥���o�5d���f'q��/>�m���v��Ux�5G_�߅7��-&��2k��eF�d5��XT�)+C�lJ*w�4=F�^ y�KmߥKS�q4Ŕ��k� �}���f��K6 ��I0�ׇ\��`���y�%c{k�@�5ѐ�P�֑�Љ8�|�Ǹ��	f��->�y�����gro(��������:�ȉ�F���k�(�T16�/VbX.�	(a��=�x��owv�f��@i��p��ǡ�Pb��7�~CD��Av�����=�]����u��n[���z)-�rQ��H�"����&�+i?�4~�0M��:v�S���s"�~p��F��+}��m�3�OO�9=[�l�ny��)��������y�3�H�h���H�༸�mm����9�j�R���d�W��J2��P�QS� }E3ɘ���F�.������3�&丅��+JVK��~��v�� ���!�U^{L�2g�~�=G�V�q''�*#���/�Tf���
s{��Oh�	��C�R�������iG^J�*Q�~�j����D������;�i�9�E�Q����8 e�2��g`p��< �(����t�l��A������<�T�qH�� �>��*�2�b���.a	�f����T��$�	V{�6T��rY�8��7��3#3v�Mnlx�	=WU�c<t*ʹ|�?�aX��o��d%���sb�x	�H6ػ�;�l�U��Ӏf�~A�7���IG�[|���`.�fa8V�bY8�@�ѩ��k�U�����p��f�	Kp�A��z��W<7l�ֆ
Ȥ<�8cూy��������Y� �5��U�L��F'�!@�m�Y��qND��GP��WfD|9��-҉ª�����N�S`����7���M��T$�S;��#>�1A��1����_E��>F���t�~ó���c��b�d'�Pz���T����Q�73V��H[�L�n�1I�����B�]!�z&��K]�r�U�T�1?w������i7���wU�'����N�#.�Ⴕ�Qi�+�)��sz��#	��!�j"�9#�^q��4
�
���V���
:WfG���ù��=�A�l���i��J��X�L�%�<�A��lAx���n�56W��VޤZ��	툳3��A�X�A�������IX� q�J���d)Ϡ��J��4.���_���wG�Ef5�s���$	����Qp����l����Y�"Këњ�3��]��F;��[�a�4�y$��[-�kq9;$F�D��܊K���)P8�LPD2ySYfE�����N�ʨ�V����R�*��چ�L-?��<�L#���LL��M�}���v��pq$���0L�)YL�[P_��捌:��������l:6���&�����n���ܱμ�QG�:z#s��`�S�%�A�m�1��9���cXe�3D#��^���B�g�}ܛ�B� ���X��%��Nm��oBWt�0�ǜ��3�kLP�lG�m)$T������<B������m���^S垷��-E���`��]HBv�%���7K�\� =1��V'x���>�XF8� ��<)Ȋ˨�e"�4�G�5�n}��o���C;d�['�TQ^r(J�ݯ�5��}��������U2��x*"�v���?���>{������b����{a��=�0�9%�利����ڤ ��q?3�����4�Bd]d9�~a���^\�OV1ܐ����ԣ�i�� �����Γ\�H#j�S�Y1pGc�d)��sZ�[�+�@��I�p��J>�?.q�,�H�Ԟ�*b!�q�n҃�g.�3L��G��P�m�n��A�g!@�C� �� �ld�W��wj���UVc�j��Pu�Q�=����P�~^6ͅ%�j���`k��m�g^x��5�z)`$n� d�D�׊k��[b:�%�=�?9�+ �T⬄$n_ə/�ل�m�  �w�_�8�k�^MVp�һ�A�R���'f���mZ���"[��Hy�݁�5��|����O�E[i�r@9��9�-���xʛ�4�ԥJ}� �?O��$�Gۅ"z�d��B �)Y6ô�U/Yna�x��.���CL�oc�V�U��Vp�"C��3���*|��єiB�<٪���f�L���I�o|�N�3@B�lR/�²�4#1�c���X���&m��,Ec����U�듙��D4��m�J��ͽ�����e���S2�+c`�l�K��e]�/_}�<�.��D4rB��ŵ^��j �CqF��~�I�0m�փ�|��3�.��������`��[)��6Q�w������F��:^\xCPK��3�Һ8́�K�����a���~�phdx�P����l|u�k��!��t�����e]�Ɇd6�aiwB}�>�����g98��]qS����Xt�6��C={=,G��mA�Ӹ�]�,V	��9>-^ɿxK����/̕ yw7��%���������y�y���O��Wg�I%B�7l�VXkN�e���[7F&�Z��M�	'��s��O��*��"��B ~/�\p�ɍn��m���cÿˠ����W�0�f	��|��� �2���+T�����y�>�4��堠�h��@GA�b����\.�ΰ��B�v���u�LQ�}��xb���W��h!�HY�䒛�L��O@"|wY��4,�q9�NZ�6�g��iT�FY#��5�>���J���>���k4����ւ!y���J��{^ciP�;G&"��1�����H�-vx���ļ>�7��_��P�I���mV���*�i�-
�{�ߢ�Q�kto��b7T��K`fzg�)0_����T\g�p�u��.�5���b�wz��M���<8�i�f1O��g'�����W$KKlk��;�FV�@���Q"3s��h�!���Lt�B>8�K)z��sJ��|���T�Hk)(,�1"i�v�K��B�KO���R8��@�1�ב��2�<��A��Z����:׷,�B�Z��PXjls�+�/���&R�stŃ���k��|�h���*	7<5�۔����#g�d[�m,�e�+-�l�no߶b=���9ᦀ���9�$lzT��H��z�.lG"E�;Cs���C)��ݭ�3��ڛa셵��P��ڪd�M}�ڒC<�����%���U�����R%a�k��X:żA�3`�
�ޕ�n+?)���0C{y��ZE���|�pNK�|���<��@�!�`dS/8����]��m0
�(�hP�̈M��)(�ؔ!�����_	sEʽ���h���Պ�'�$�!k�eU�u�������q�\+�ͤ��k\��G����A��?%�����R��wWW^)4�4N��a�$/��5O%�ӝ��3^��{��� >Ư��vţ�h�\%e�=�B'��� k
VX?(��]���-���%�u��ce�
��Ps�Nln��_u\4_����XY8�E×��.�,�n0a3�X���@�#� ∥�Igc#�P9�1�[���ՀWV��}TTŹp9�a
���w��xf�Ӈ����I��sb��<�F��xz*��?ژ�z��5��i뾻�)i�5LI;����㎻GA�(�S�t������yk�$�ҍ���)�_𫄃��q����TIɨ���/9�Zb������&<-�B�v��n�9�ޖ7��j-8{��$u���b8����ԯ���.��o���t? �/m�e,��$��@�cW���wdh]�,���p�yUr��>WO"g�0]��'�Sa�ɿEr��}
�5`���J���Kb���/\E0)�~<1C)�t)�6�iH��+^�
 �i��Q�P�(r88���G�U���,�Q��A���s]Wk�I�Ϸ��e)
��;F��/����Y~���<�Hy�A��$��&(���Ni)��F[�}�1��qmo�4���7ep�T��R�|%��I:���QZ�<f��M�3RR�,���]�J���g�t7�����]�X:)����X>f�M�}��W���=s����_��>N��+W��c�V&od�G�T%�n���������5_����萓�1��YRϤ��Rq�R� &P�g�a5�#��F7g˙3� ԚZSs�����2Q��uxnaۢ,��DAuR�����T���%����Q���z�@�:�ߕ@��1�b8һ����� {[G=Eg Dt���E�G�E��X������AP�#��5�݂��13R-⫁-���OTD�����in`jZU�����Y;(`�����4����R(�i���+̗`���7;��ގ���)	WaB��:W��21s^d_������#@�l/Q�b7������c;(�x����}�Z39�1c��l4Y����%���D���:Q�x������m�.ڈr��@�b��Ba�u����Є��s�?�Ӻb�*Y�*a�L 5>��ng�u�����5%X��a�Hk�ƘuI�.�h,�����!�-w�^�o)V�?�Vxef7��O�q�[��Ed��c��~K� �;��`E����"�.��� ��-|T	4�h��=.B��=�dTx�d	D��;f�wV��%Q�����
Ȼ������nV�9"e��*~��?,p��I7�<��#����L<�@g={᝹��C��H��3���b�m L!�XH=	��?n�h�6ԓ�',L���R�?j@������h�	N0lm0�<���-��cP=X%Q�J_	45���?��>� NLG*.f�_!{��|�,]a9�r"��Z�?2��ZZ�{&m���B�����E�fŜ��X������+KTf��>s1���p�2@�]�e�c(�Ɋc�3�<�B���Tڌ��HЂ%�Y�{El�ASY?T�I&WxAW��b<	��T�Æ�o䅱�uV�>�� g�ӔP����"�8��N�2��G9|�Ю��X��"��e�ʁn��#�ֺMW��Xu=��<@�|�+����?�7^?r�gj���#k
�?Ի���A�TY@���`�6����@���u�� ��_c���c���R���x��R���l���P���WGj���������-16��i)P}�.��`X �N�\��u/MF�Y����s~�s,C�*�gi��J��@��vo�-�wlx� :BD����j�3�zeouEܑy<�O��^��~����Ձ�����fR��M��h*Z�~�e5���V�/�P+�R C`������i'4[���}ܭ�*¯Q�*��HJ�7�]( 4�{�,��fԺ��Q玘sW�����!���G`�I�R>��5���)MeR�H���;�M�ED�s��7�]GM7˅U��>�o�����rTX�Gj�n�d���s�,�]F��/�:_H5�����S�P%$~�K[0i��ƢpZ6�B���!�����?.A�K\�5wbSYX��w�]�~X�ύ���,��4����NU��?;����J(��c\I�E�*}�wF����Hfs� �L xmO�s�e+$��r⡦�
�@H}: J%�����o��w��w�f!z��y��	�fV�00��,�p�E� D���!,�;v^���c�w���X��7�+Z.�gT����
�p�0s:�A�`EZ��&*%0����#EYz��^4��g�x����Ƕ�(�R�ǟ��:Ʋg��b��Q_�k�)�lF��f���&N+@�y����t$O��-��Ҵ}�.��?YchZ�+.9��AO�YR���dF��l5<7���z��"����M�;���1�9nCo��?49JL��H�\#�i*ѣf@U{�b������)�����U�K�J�����J<�`�Q#����@�zx�`�� ]v���;鞈o��aK%�;���[�!x!�
��Q�,+F+:O	���.2��u� �N,ݍ�,$!\��mJ�B�p^1��;Bd�mM����r���A��Ϻ@`!胪W��
&��PB�;M�>�?l`��p��P��C,4�n�,I��/F�r�u��;�Ej�}��x�J@��[܉�g��_,.��&�A��s8{8@��T;^��R���>��C��%P���4w_��zwZ<� ��\�29���ND�ŕw^�5�RSAG�N�@�����ⶽ� i�Պ��t���f}��|	|�p]�ʞE+����+�����a�E�S��j����-�B]^ѢQB"�U�*�"�5Y�_�
rp1���V΂P�ߵ���)HAU?)�v�l��P�YF����ؼP���[�'�Bl����/>�50b�;�f�n�b��
��j(����#��{<q�_���y�w�p����+�������@����h'b�'t���N��v��"�ʎ�ܝ�L�s8����������I�X������g�+���2�S�f���IYVڗ_��ݞY�y5�N��~��N��4`��8�TD�����T�Aj��_��0�@�A��`��њS�=Se&qt�Μ$�{��LSN��K�[Mt�����9�׎�����]omN ����سYB��F�uiU"k�ʻ���������+U������8���B���ċ�y��.�F�m�����ҕ���K���v�F\=	tǙ�oO+.l�N2��唞��	�ib�!T ���y��sĭ��r�C,O��8�z��|RB6��4^Q��e����/��I7��3���ʞrc_K=��V�s9���kKRE��<Ͻ`�-4A�Hv�t��w!1q�Ω'H=�^�[��-�o2�vG�V�s�����V(�e�\�|����p!��ȋ(�� -oſ�H��С5�Ȏ�W����2����t�)Ԟ��sԖWA�����[ ���6�K��f2�d����4�5��ス�����ߴ��&y��/Ֆ��O�}�Q���r���0G�6 垐d7S/���Z?I�E?½?�^����t�j;�"�����Thʯ,t��'�u!��1ٴ�w���>�����Gz����:m��..�o�� ��
-���[�~��C����Q�^�ji̓�I��O��z)�$oQ��t��'�u��R�2c��ym�I�;@F���`��@�E/���P��{� �x#�݈tNRx�?��$6�Lrg�X�`�&pG��+�1k=�:��e:��-�P� �$��Tfb��z��a�pkܦ8ƍhI�S�\����*]��@7��-?B�ni�G!��`d�p���"����0��b��,��"I`}P��&���ո�TC����C�Mv�U1��H����J��{b��%S/e�΁�!I���b��JS͢G_G���n���t��4�;A�.ae�%�ߤ��4_� �Ȱp��&�������2�0�"9�!�J��e���$���}���a��'��ǥ�����˕x[Cz6)�����r��,��Xd�\P����ΚڈL�<�C�F�򙹃l���30֓6��0];�����l��a%ۚ(�zK��B�l|�$�I����ξ�x��ԝ��IS��0ȥ76ev�dio�Ԙ�&�X_N�5���,M���� dw��?j�{�S�
/��X<����� XS�'i��?�RaA��C ��~6���$(77��I Z#Nq�[�eh�	C'y�"B1��<}�@�7G8�|D��^:�X)ꨳ�ddS�F����W���U�b��t��KG�Ԩ;P�F֔�/�\k�tt���*l�?wfd8>�Hb�>���dߎ�I�?wZ�|z�<*�3j��g�O8�s����m~R�7n��`;P^/'a%�V}b'9"�З㩂<qť5�q�ʁ^2s9e���TYn��G��$P�@9!}��K���yה���cŀ��/(���r�:�&(ҒL ��"b9�Dώ�M|W4�e�+�Jh���܂ �p���sg7�l��D���DmڔD��\��)������ȇ�s`#���]��݃�2��ui���Ď$T1r�iof�X�ɑ�!�j��?��:p˺oJm���T�)�n�4 q��j;�����h�	�Ě����^�h�uZJ�װ}�~�|���7�P�PAf�%��7��fL^�X|��D���i�67�Ky���,�ߑ;Y�D!����3�x)����Z9o
�$n�Ը����m-S�i������o��0\>�+���"�~Fo|b��(�CG�� �5I��dZU�V��E�{��x�_�ѝ	�'R;Q���x99�
^�*{�Xͪ�y�*"Ќ�NG�<�Qt)
��Lu-,b6'"Qu��;T<0��/�P:/1`�>�)���3�W�a4.&G̚��5��M�)��
��	|c��؃�۶�7��`����I~l��h�恽Ƞ��_�����\�kB5��dc���	l�s�����+(�mmma01yŢ�iՋ� �NZ����(k{�T�1��Y���g]L���͗��3{�Gg��~��k���Ǿ鵒�J���*���Y��ί�X�=�E=�Uo�#��b�/��D��]XBC�f�;��p�=E5˸�B����I�ѹZV(4��46@���b�������2��~5(�.�N�E��k*�A<��ru<����X��a��߷��T~i�Xb_�#*�����{7P�<V*��0�B���j�`4]�I��r��Fsk�4߈����"D�!T��1>k����u�'B�nr��2kBX?�2�؎=?��m��#Ի��d�٧�1P�m9�@�,�����6�Q ���	�JB�ͯZR�������S�"���܈eɏ6/�xf��2�ݷME�L6���ͨ�,Wl�*���a����t����,y���#�.9�k0@J7(01?�1�cd��y�*���fu�b�<��/.?M���_0�|��K2 ]�.���cR�qY�:�Zh�/�'v�`��� �[Fꞗ�*9goGePͻh�H����~݊)�]D�5!�|���
ҰU��9���Y��E|8��Ů�`(M"�Eza��H�x��g��X��}A���^o��vC۶�Ms�O�ߵU����S�8�M�dn�@DV��Jn�6��ax'l�j;�󜨾�@O@Uk���E���Y�id�%e3ܷ�Ƽ�W�L
^ d��b[�M 8��&0VQjt%ѣ�b?�0���pO�t(G|����W��20p4��D���+�	�a5�`�V�=5k�k��Nq'䔹8�[w�(�����/�ck�!S)�`�0��+�Q��YR6v��[B���ư�a�'�䋷']_Ţ�v���,�|�cB:�7����!�D���_i�h���+S�;��՚U��|q/�{��.54�q���lS�i��נ-�T�_��k��Ҭ���D\?.���X��w ����g���.?��)	��1����V�*\����v�eA�<2�1r�DI3�XT����7�_~8���4��7@����vzOۄR:P�mUépoUYxe��3�5�<�16I��Z�0h���f�I���$��E���}iUZ0���R��V_�����tKB�_��10l�$n�� ��-�X�خ%B)+k�����6�h�'�C�U�Qa�J�w��TjY�K\}Rr�ö{4�A2�2����Y�^o�\���+� q?�%��q>��Wk���R�q�6��w�7wObm��� ՗�1CO�\Gj��[bT̾s0˱x���7�H:�-�=���;l��]���,(��8o�5nDl�T�j1����`���}<oX�TYCK�"Hg'�h�i+W�ȴN�� F|�d��,��çl��������I�Z�f8׾��Pd[z���0�7r��5i���p<��s���ߩ$-����1�Z�_7-��˟�I/���ҚX���i28;6n��;PL��aq��5.��g�}�WJڋ[y@��J�l�`���b�����ǢdR�Fq��E�|ȳ��n�b� ��\�u���ɪ�*-	���c!��k6ur�>t�i��N�����h4@�{Y6V�7JȰ��-�f3��+KM� G����k��%�B9!�9��st1��`�{�Gnu��v�?�V�� �q�M%0�Ŕ�{�g��2�~��Ia^�j��U��9�w��f�u��˨��Q�CBY/�>6�l�CK�<]�1�eP��p�xh5�<�r����f���^ɥ��_lI	;��� ��>4��|�9��y�Hӄ1�Z0Ǟ���Z!����Sܙ5_+6����{K	�y2O��j��D?^)|�1�"�nꯤ��vo�(h�����LQ�=`��|�Γ5�d+�u���0`|�/���ϟ�\�bA���~��b����C�cJ�/�ݮ��Kz��k]�^�o�C�x�(�Sxcs��D�yޕ�:��5>~di�#�M�
��j�����-���I�"�a�&5�"1���{���퉳�?��1��<>�`�p���8�5El���5�{�,nV����^G��L*d�<���%��AvQሣ2��zd�Q(�m��x����H�H�q$�1���/�V��NP�W��\Bϕ4�X��(6��wk�y��jO��P8��f������5,���-eCx��]kZZ� ��A�᪩��I}�&�Y;֣�b���[�(y�3F_~f�Ѩ���/�1(�kl��FD'�XQ�ueҫ��\�n�{:fZ�{��W����`�*�6�j�f�t}�,����f��o��¬�ʹ4N^�j�_��� �\�Q�a�B�i�9�`�MFF��ShE�^u,v8˱� �<��+�!�𧧞�=-��SP���L�|}Jh�
���n��x���7ہ��A�XFAS��I�
D��7�V3�'(_��N]��؇�1h�|���	T�X�v�+�	��kńܲ�n(Uժhu������j����8{٨(�z�sx��r%��Υq���n%��P�g4�Go�)����>?BN�gi>�h��):�t�D�*b�J�9��"�9��`Ȑ�P�G	��HqcI���M�����-�[j{"Lvj��������HV4zZp����$�G�[�4^�� ����OH�z:�52�*ׄ��e^��L�Rv�!�aM�r�+��f.�ws�&y�LCM�f`���˸��'ύ2­�;fH
�M�/xV��t+{���!��F�B�@��p,�x�s���vd{޾z�v	j���+L�N�C�(�a�����x�0Mڂ��Ɠ+�*#R��I�,���v���7Ķ�?Q��>�2R�+��U;�(`Ue%�D����1��y��ླྀ�1�Ci+*d"xR����:�tC�=�=��Eً�_�G�$�RN��12��$0������+m�C�	-��Zg<%,�']!�I��!X����m�_��JJ��Aؘ�树�"�۪K�jH#o��'B]޸G)E�nN]�����C�����T�' �a �s�+�����4��XChh�����q���)�������#.�DtQ}��gHl�l��d�Í,hJ|���2R�FbM���u��a;@g�	D�Y�;�1���]�ŹwmX/ʈDg�^�{ɔ�S=���0���)��JB����?�t�W� �����񆶁��#ÿ�MWIr��K�g	ɴ�"o~���N�����jڿ'e�1XP�K�f���`��1�j������K�D:[���%eh���{`+[���ȑ�W�n�X�p��A�4_�V�����[��mV���g�n��ܷ��-H��>����[W�g�xٺuh�R&롷���?V��_=���7�c�I8���zo�5?��d))�$=�1c%1�9�Y��VЌzg�H��vg�*$�'�Q���a����q��i��U�ъ���X��MmR�8{բ����I����I%FQd���Ԗ+���P���':!��T ��%<�.d������T�:W��]#���/�56�,�
��E��7�~���4��G�C�,���B���@͵UV@��u��Dn|����';.H]B�٭;O��&\����
ѧ[�e{�utK$��r�s9��C����&j�K�3 o�Y�,v�|cC�8�Sf�q��awd�������:2�X�fq���%7�_�L�׃�Yɶ�O[�0�ᐻ#���Xvґ��gi�ۏ���:®��E�ˎ��)��;���*���*ׄ�����	���%�3ÏlجY�_Á�����e~#�4�X�;r<ָԺ��S5�U����i�6?&u�cdB�@n�����ɫ٨�����!��FSPa��V������\ʹ�ޥz��B����'<;ߢC���#�Y.l瑑àn%��-��Ȳ��;�:�*�ĉ[���e���l�P2z�Y���D�1���Sx�{�j�ivѯ�&����#B���Q�_CM�6D둊��3�@�H36T+�+�Ju_q�"�M��J;��p����������+2�'E>|0A&NG�0Z�t����}O�E �I�������`'�\�h�v�AL����Pd��4zP�k��\�K���dPw�!~N�1_ye�mz��`��H	�x��'��G"��~lO����N��7��^��^F��	����w�`m7� Ą ���A��}��-}��勯E��(�)������_��w4,ɝ���B\_ 	B:��T#�!�"l��
�~7�N�"!���&��Y�^~jH��`:���$�r�o����?�p�A���
{u8S��!�@�|�Q�=I�R�`�=��pVr4�Y��뭺�w [���5���Fw�#����wR�P?~[��lfk�A��+���fp%׆�"��
Ǩ���K6�y��٧�_r�JYkܥ!U��;ʍݳ�L��ǽ�<��xa��3>g.Z�VUK����w�ٞm9� :���k	�]�k�.�\��V hW���Ϝ4n}a֪���2Or�)	g�룒�[�_����֒���}�H*��j&��5�mL9��x��_�\ҽ���L�؜m�D�.����G`Q��!v���-n�aY[f'�S�]��m��	����zc�sN��E��\�z�rQ�p���L���} Ţ���'�E�ߎ���e� �����0�+�%$�� \m�ث��*�4���v����i����X�z����ƨ�eeq����j�-gcE�$F�_��-�ū����K�e�3G]�U�7{_�0;L6�'�V�^��T"7�Y��KU�W�@eBӓ�`��I�$�Z�_��oq���k���XX��7PC����Z%��+�B�W��H�1 �'��B���� �_ga4򖌂+���-���'�ώBf�Ś_V�=����� 8�Mkfe�n� 3	��Ex.U��3	T����po#E��Z�"�秛͡CnP�|�R{�J��>�q!�4���y�C�M+�*�<oU�f����'�:���������})Гڡ��|i3�mYߺ�����d��Aa%����J��j���3�T���{�ҡQƧј�d���y}�����2F�$�SYY����1���`��"���žk^?�+���w%���|�!�=�d�jy�W�Z�������!���ϯ��1�)�-2���
_5]�̠hqVc�-�݆gI6Z4~#����T"�XM�Ֆ�O��}��
x?��&���[�s\�`��4�T\w��wY/�@�'{�v��L��I�U6��g�<CN]��)�)Gل��#�*�� $P���O��An�v�"�M����d�獑0x�RZU_Rc���d��'��Jfn�S���t̬�"n�,Qa���Y�p����(U�6�0�QR��0�3�Y�& !�����w��k���%�5a��-����^x(�K�%qhrA*.��rS�l���ѫh�*��1ڞ�p$ ihJ������x�r;L�Z���L��h�P߭�O;�WH�y��d��;f*�c�����ӎ
M��k��]xSa�[M*�\Ѓ<�N^g��4!+a��!~�h,�_��y�\�̪�'81�.�+�XW��*'��-' %"1:�V�&%��(��A=Q�BQ�Q���H��r�ڙB�,j�2��=K�7�1��z��.!v�uh�\ac8ƳՇb����� �Hp��2t��F�h�+漦���-��\t-��5o�y��ά����:ƅ��J@��{���?`cha���XZ�j��A���*21��x�У��k5��J�蚠B��Q�\A�:�k}�P��
r�=���g2k�v�1݃t;e���0�t��3�;]���
�ʚ�]&�r݂ٮ�8��g9�s̬ǳ
wT_���βTkh���M
<�v����,r��:ۀW��#�k��:|&�njL�rG���ݙ�/�e_C���k9�'�RJ���x��[t��A�B�c����ӫ��n�I���3�,��"��-�uU����pF�O	q���˾�f�xkCT���>o& Һs��q��Z�f���?z�o�Z��G	�����D���z�j�Wi]�G�������D�hI�8�$�=�G]x�x��:(��IА��ń�xe��8����BWI�'F���~?!�u]p=��X?���ڈ�i��\ܝ�✺�*��D����i.K/q4*�w����}��+e5��Q�w$�n�����M��q����x��s���ӳrU=$kM
VQ.F�V�c���q�Q�5�uG�RǑ�9�I�*��6[i����)��o��ߤ$��t��h�eS�1X]z��R0�7k�響�7��4��()|PKW��U�=w�e.K��i6���}�����x����j�ǵ� �γER�b�tX�a�/�����wvU��B0V�/Wnt(�S��$	�=A~�Z���g��e����--At_���v��;��'wI�C����f�d7��������C��SA�K`�\�&��0`��gCSO+9io ���Eo�&��E�P�ep��1�$�aS�a9Qp��r˦�w���ׅ3�s�?�$��q(��1^��9�Z��+'yxX�c�ܝC����U��x���u�='�@bd������H�H"��W0Pc�r��Э��.W/V�����!3khp!��{1D	��b�{s�p[Kr����)'	=�z;��"ׅu�LKevA�����=��Pk9Т:~� ��b��	��a���o�'�D>��"�@u�)�}����";��-ϊmtl�šE��mY01p�GeT~Fݸ��٫�~���s�v�-�Y�w��o{S�(�#��M5][�wꔅ���!]��ճ�Ň�`ZI�����纻��@\~�a�{�H(�rX��Y�T�y�="�͛`�Ca�#x��8uy&�n�_�����z�B��$���+ۿ?Ë���˭�.�I�+��_>��x��&:,F �:���HZ%V����B�6A$���ߢ��sDj{4H��:�Z68��X�]�H����������7*����9G}Q֑eetIl����Ylb����nz�y�_��ʄ�Uܫѹ8��[���Z7'-�(Ox�q�ᑡ�H(�w��;�c���z��&c6*5��L��q�ւ�(��u���Gf}a��Z���d���@�x�0X���&|�*��9� ����Q7�Q�c�0��Ԓ��#ΓB�8�����8�=�
C{���� a��H9E/�n�w�s��M��� �z8�.��	 H)�j�Z��݋|s�}����|���,�]r����iX���`�Z*����a:�cR��)E�o� v4�8�r����#$��l� ��Y@5.�HT�2�$=w�2��ޚ��u��T�KA�3:��<h�It�n�����|�cl�i�J�k��2�ѷw܃3^)yC��S��dkyn�����6��cb5/#��eU51�ş�Rc�{O�*$�aÊ��"��t��|��گ�IW~�E����UaH�1& ��|P�zy?9LV5W#RZHSE���_�����[���'�iϱ	^��1u G�H����/�ބ�LJ��b+�����aF���Fg�S���x~�X�\C��ߤ�#0RdSE����T&����T��Ţ�%$)����C2�+Q�i~�1�3T��N���� a���qO�s�Cvz1� �^g�`p����;+�Bt���\ �B�]k�#�,B�Q�So!�KRL��L����n�����"X���:�ƈ+I@�b.��+��p@E����jL�R��E�((D_���/���l:�xą�-0z�������xV�q-�']���gT0�Ύ�Ơu�ҙ&�M(
���.�o�`���p�&�mC?R1蘆���� �SC	4N�`�@�6�Y�� kv�pR����LvX�<�Mㄤ�4���}�#�ÂG��y�Q��4i�7����s�I��%��[�jh\��P�J��ſM�/R[�=]��&��,���. +��׊�
��˳�K~��)��NJYX���(>Rdq�P?2���fl�;�rF[|��iWGO��M(�Y��_R�7�a��*\�-�2��&�
������z)'�E��H�%��v�˚�tNO���{��m�����h�<�וzF9�G�,���6Dc�=G�R��5/�(�O{�������a<'e�%>%3��xNg�d�50
C�d�w�^�P�@ßB*,��k�@��v��ٸHB{J���eW�S]a�j�" �Mk�]*�����R+^�yNt�%�2���x����Y(	����� �>�ɭ�Y�؎��f�s�_ӗ��37�eF���̖v6�'���֗��J�X~����=�8-��~%K�h� k���4��w�S4]^�V�NR�m7�|�U�bh�3$�{x������Ȯ�;/���1�x�p��14c�/<��:�p91��ȫ3!Jc�A��<��Wc	*��N�.4�>��e�*%�1+O���i�$m��5]?�9���3��#Dv�Sb���]a��N��Y$�oS47d�-HS�Ttb�y,�bgi�(�F0faA�uݔ���{f���S�<�y#�F���X��8 >�Q�m!K����)|R���ʉ�2��o�I ��,���v�FN�ǆTm�a*K Ƿ� 6����2�`F�o���D�M��;C�y".dl������ク�Os��v�ҔtP`֌L���$�2;��z(�qz�@���/��:�Wܛ=s*������15�(���p��-d1��̦�����KqeW���~:#�,?������Aa_���§;��ד������}U0�� ���c,v/��ٱ�Y,0�+%��/�2��|�[��c���)�`M-wF	��a���E�5�5�����"z��RRWGa���zOYIv�9Cʩ�R�f;�S�-T��ܒ�cq����#6H��-�d����/�B�P�"�07�>6�ې��F����1E�����A��S��6��C��GQ��
R%�E˂>����Cs#�"k,��E^���M#ĸ�(3uv�d�C����iv���^K�W�q��yJ��Z[o��C�jvo%��>?� �w�}�&�� � !8�il�IVf��Y5xI��%-5	>(�Sz�Ky�ȗ������X��M�U9W�� -�[q�U�v��"��9[�(�#(����.G��Ky�r��z#�( �p���n�,�om�}���ȧ��̘$JEZ�W��/��H�{�LS��|��D��+BT�y?�;�a�1�m!��4��$�PB��^@�v����{�Px�����>��bk�9�\kst�MUcs��Ip7���˦Dh#2y^-~�:!�����?]$�YRD���������e&y8���GCa��RN� \3	�<�Z$��ا�t�����d`�{��^cyM�Y`Q��$^veW��M��nZ�"|��I�r���J@=n��td̟���D��qc���q7TƋ�,0N!��9��17V���D�+볉ʈu�+�� W�M)��мh!b��Y�eL<��t�D���G����)+�O�v�䮝�y�9���qw��|�f�/��1�卓؇��~�˷�֓�{!&M�#)�p��<:yF�T��S�����fE�p�	��+E��.L�iG�G���n�:�b�_;钙���j���Tu}>���9�1� ӝ�U���{wAm-�m`�����L�2`>\�#Jv^�� aS���x�%�����ί��L�k����z��c�4��ׁ8��v=<�UF��.���Br�u�Rۑ���s;���M�==����:3K���0��ӼPsi,k�Q�(�u��
�L�i�<�uc���l�{B�u�&�����7���uX\I�r�X �;�(XL�i��']Zj=��S�`�|�ګE��%�ӳ�� ox6T�c�}O����58vYY7��PD�L �-����u��A��֐���fVh�@⊦�[C��NZ3�X�vL�X,ċ�li8b��a������0��ҫM�5��N��",��5�5
���#��l#@��F��mM����r�޳~��/��Ra�������D�N���! !⌖ϰNJjv�=H�z��+���`Y�K��W��|DF@Ƭq�f v�o����AV��\��*�a��fl0h�$<��u��򁾬E����� �3��x�mpwǐY.��JR�	����]����e�	�襖Ӈ�*=��g�&����oT��Av8��\"�w��a(��`����O�3��pk�Km8+��Ӎ7 ~f�c�906���T4�k�r?~T+B�䧩eTR���"�vrL_!�Ǿ9�13nE�����i�&�3(�X�hY�sǔ��'F1�E�S���=����3F=���9	�e�m���v��
������x��#<�1�ᲥG�;R���Z@G�<?֧!(ټ��a+�咨s�B����Ƽϗ�b����X^�%id�%�j�>�V0[i;#��g�eMZq�^��
�l������c��|ɼ�b4!F�#��C�Q`���ֽ����^��}9��^���e�	�:\�m����	��Գ|���a	�J���{����*(�`�t*�s�#��M?�j��a~������pb���;�4�!�^|�@��9M�-�*[��#*��n�I������i���,�j�М>D��j��7�GO�9"9>ɬJĐ�Bh#��oC��nο���*�K��4s�oB�nJ:�G�o��
�Ǣ�d����>Y�a�ϛ�U�7)L�����ͽ�V�+�&��Y���d����\��u�T�4,%8�{l��~ԣ�V��`�)��RMv	��^^�O$�B(�1n��)vn�M>eR9�ꀀf˫_����J���8A�w�CrS���ʷ�����od��4+Y��n�t8���QںL]�D_"����ot���x@��߆f�My��&�*�{�<w�C>w�p����|F)�xE��RɌW�u����̠�(F��ڏĪAi��h����Ǻ�L���
z�l8B�ߒ0��Ȅ�ĕˣ㖹��}��NzB��Z�=�2�JW���5~:��^h�C	m�[�_훔G��+bo���K��J�y�tUk��7_?�0�#�)h �po�>u:s4T�"?4}���:YQx�Y�v��3����SEo��G�Ϗ ��ȿ���ѫ0 �^V;�6�`&()Aȅ�6^�NHfX ?YC?^���ms�L��$�1���`$��!��2��Y<�j��>�M�nS�@��P F�a�`�m����I~����W6E�g����>��Ū��
��qȠ�y���7;<ٝӔ�J�'k��8�Ot�C��d���_�$��>Ԟ��9^��ʡg�4�����B��'�����૓	�%sإ�hbR���
Z3�J�-m֩57=�P�y�i���Jl����]�Rr����"A�Hu.�%ǡ��`� �/v�pA�~���)�&�����mXeۣ��'}
���L�,.a�{Kk�HV����^����L�nD�AJ�^#u�e�c5�+�U��~C"�2�e[��/�{�f�$.�̰��wg��`k>şoV�Q�ÿ��ߟ��yI�!�X���w2O-�;k����W��<���(��v�mlx�)NW��:"yi�{'��y9�f��AO{�����lj��J��p�T����w{@1Br4��*���:�d�ͯV�M�L���ƞ8�|���cWɽA�:�	�׾%1������r�� |�J�.�A��iެ��(fI�V�Sè̶#]�#����r7eb�Nܒ3���I|D��L���u���??��ޫ���������Ӫ$�z��rhP�D�7�??Z�mYw���~^TF_e�/�������z���ډJy\�nA�93Y��f��,C��nfܵ'��WZw{{�X<��i-[E�rI�zD4��gU.�.VU&�_E[�I�*�&�Lw�*�%x�Ma�v�+ީ����탥����f�q%ǀ(o"t�֚b�����ܸ0�"�M�<~���UA1pF�9��KF���,�#)�{��w��:��6��#Z(UD+�<{ob�	���Y���YY�Wow/�y�>Nf�2��,pnb�޽=��o�B�
�����2��l��f�q,^oBMBp�X)+�8��"b_B0Q��[o24'Jk�*`�1GF�t��ݽ��X_5�|�������� �pA|�X�T�H�����e�	�dhO�7���'��9�ѺC#��Vձu4��	�����vug⍒۴1�z�D�9]�e�8��5"}��!��"���D���F.1��kb6�v�����*RI�,K�tW5XVU���T��q�|+,\v����"��gq��nG���(�ʲ�ަ��p����80������8V�'Τ;`���G��^�A����{����0[Sy�z�%#�\��Z��-9,Ec��P��MY>"W�󜮩՗��=[,Y����#ⱃ�,�&L�3�1
�9��x�_x�0��Oq�E|�"{�m��z�V/�ş`.��A]V���r�L��#S���v(ԥL�d�c��I��H�r��dݒ��J�.|p�����+NY<�τ�hN�RH�T~�ѽD沪��7�}K����.9��<���pD�><�L_r���k�_.h5�ڂ�x%�����E*�|##�=�b�0_ߛ'��l��exG�ڳvPK�	����WP@�q2	Ə�[���h3t] B�B�tθ�[�"�l�!�F�/'�³
8�% "���"Ս}��hg�\����s]ϴ����T��\KK�FЪ����5��~��x����U,ΆJ�;�):�4n����xY4`6��/��Ve?���%1h
շ�~2y��'RȂɨ�3�P$i�ޞ���f|���&�v'�{����x�w�1sm�W ,��0.\�3����9!�~CI��$��se�&��4�ނ����L��GK���(�R�_	Oh
�X3|]�j�/2�Q��=���MV�����Ҷ���Fw;��2S�v�ʈ�eb�v{�]\XSDT\�e��;F�I vA�Ru�`���V�z4mN�P�yT��WY�WگJ]
��,������D����~!g���a3��ܝ�*��|�M=�� (����Ǚ���z6o��i�3��=�(옰�;R�a�b v�{\���k7�\WI�i'�	�+�+����1��;-�#��I��	 �@B���|�c��F= #�|�}׾�Y ��՟H�KQonc'0��tW
M���a:8��1~�!B�>#W�ݷ���	��nl��^XC=�O_;��E���[�����P�Ŧ$�k:�/ΐxDҮ��SC-\pYm��D�]��c�DI���5�r��+�������i�ҲY����@�{ޝ=�����x�墠B�!D>PaX?����}B5}�w}C;��&5��$����H�-y��%EF7��Jl-�#a^�����}�t��B�H<�_������.$e���̼���պ3T�-:���F+.>�}�n�E�p)��
F(�	c�Qi@pѳO"f(�ٜ��$�>ݤ+�4()ý����AP=����ܪw�VA�qs����A�l�ev�g�I�MSp���h�齞�SD���P�O���y�OyR�;��]z���W�F(7��h��|�h/s
��c���c�~hЏ�-h�T
C6(ǌ�Ҁ&�普�;��O��� \�\��L�i�L&�\����i&��\���D؛�(�kk&�Wp�g�I1)QvI4m
Z��uT�d���,�u+���&.:�Y��<07L�G�_��"���}�������p�0#��%U�;>S�Y,|c��='�l���X����,Py��%O�yD^Y��7��)��.�.�٨ �6D����7���5o��h��'���"�'���|g[�v��'ڀ[b:�嗈y)�������R����{c��	7���|�U��S����L�ҙ2�����$q���^><A�>���)����3�|j��WÄvAܱ�T��$>K/\�]����k��X຾�Ɍ��s��e�d!�m�DY��Y�O�2��0W-��#H[��*��j3��� )�]��O���q�:ۢ�����
{	c��Wy��m���cZj��)d¬��_m =ŀ��)����4)砇�^����)_9��y'z�����~53�&�?K dO	�8�ִm(~�h!y��.?4K���no���:T�!T�@~!�Z�DC6�WI�@��9��Y:�"7��T�
?(B�n��I/�'�V���R��im	��lb��>��^AmO��99���4��2���KFQ��{&���9�^Q���~��Jn��aʶ�=�c�>ˍCa�Pz��`�xo85 ��|�C"lNu��[a'�	S�5'���;�=K��i�o�{f��h�J0T8*K5�|i���UM��j����z��)x�%"4�ŽԐ ^�;5���$D��m<����e-��)5Ǎ��q}���4A-e�{��{\9�~����rs�Y��&�n	j �"��>�$�qƥx m��6���-l��Rd%�._\�1�l�?�h���oXK�X<W��*�x�����N�8�e�:\Eϗ��P��`n��A�k�&��"̷�����_g*���QK@������� �AD:^=��q: um�h��/>���!��՟b��䏔�тz�o,{�s�	3�W�b����Z;eCe�Q��	�&�Nd�������@�Y}�2�F�0�-3G��k7���3P]S�����=	o��>�o�'�'�oO�r���ٽ΍�����)'���b�l��'���a ��D=�1^Ȟ\��;�\��L����e���ƅ˃53����ʗ|�9_x��5RPR^@ho�g��f�Rc��+^�ݸ�c���{ɵ"F�Z)�%"�*�UPz5�g�@t4��{_��MOS��We�wE�:���\kx�]���r������n���x	�����3�W_��.���@[j���j�E�u���'3U�T*�E;a-���{X���aq��~��31 �em׋[c��3�>l<Eh�
TDb�%�Z�h���&N�aD%�x��ou8\3!8{���[�j���ز���X��@��ħ�6��I���	:��:U�g�a=��x�=� F�C�+����S)��߈�#V�w$	[9�m�E=��S����g��j����b	��|���������Ê�ħ�%�*r�5p&�4V#�?e��}�{�z6��m2j��,N�Y�VnO����3<b��ZSn_ב�'M�!c�W����%͆ ���k�C#����NoãI���J� �����j lO~��^'�����pUf�j��������k7�Z#t��{�l`S���Aų|z��|�8� ���q�s���M �ҹ??kF���xw�0�ic�nLၜU/;�`<Ecn?�m��3�x����Y����\8�p�|e�4kS�c��|������ض�X�6�����8R����w�X��Zb�h�@l�lC���M���c���Sc�,/탖�N��<�=#P|b/z�עrA�t�Ǘ�0v��4�/|p�M�T{����uv�$��(6S`�zم>����mT{\���Y����<r�C{��1�Wu'=xfH���8*��:ZG��*?�=[vo1x��s��F���O���Oe	Y�J��^��4i�����)=�Գ�ң�qG�΍4�|`�J}gt�
۽"!���1䬡��0�0y��٭1�ڛ�S u�YwJ8>���\s@b�/�R`g�D��v�[C�ֱ?��n��+�pˏ[���H(��ńB���t�d�����hx2�=��Fv��.�����O��4����8�D��\�?�]� f�KY�$Ƶ�-,��(�Ϸ|�H|X��ۈnc�&r]������H��~�5�/R|��D�X���E⟻�"U1�D�\ݼ�kK� U7�/���KH���i�"نZ(�tn�V�0� �ԕ̐�nYm�7cf1H=���d1��^�������IG+�\�O�E1�K�M��� �H���HV���+�XI�U�Y��2��{�oV~vO)t�����c=|�y��u�S�)Wo��YY�L�x+&u�w�a�{�vR��zq�'<M��	K?�:s2H����z8N��zx`q5�u˨���TV�� ����E�S��T���z�xF�1&`���l���6�)�9����0�K ��?�׮#]$��v���,8`8,���<H��'�QnV(MVN�1`�A�[��	V�S��I-Ա�,q��.�rK�+VҴr|��Q��B=�s�n��ckl���K���ф[���w,�~|�~R��:�&��|+7��l������f�Ή���b no{!�Os�����5���ֿկL����;rEsb�eVc1���:�p���ldIvA2Of�O�����>��|'���� �ù�{�������Gw��u�5�yYs��p��V4���4
<G�\J�.���d����9r3X~�<~��ֆ٠���}��SԳX׌�qIVHT�'V�\̻�0��@�V��^=Ծ��Z���pyW�L�>Bq���J:ɵ� .9[8"��e�HU-ߚ]���S���+!k_�(kQ���ub2�*�6��|o:�E ���� f.88,2�Kr�:�]�N��/.�PWe�G��"+��%��&U����xq��Vݔ�8�d}Q5��f�&X�D(��� 	��#�C�F� :7G��L�i3`c!1V&�@0̓��u���q��n�a�י�ܗ{�>d/tC�2������¤��\�k�sP��2h�
dzׁ���V�����#�C�~�WIx�c<��#�T��7G)i��M%�xHYKN,+�	��vv��?��qT������o��B!�fm5Q�
�F�'�4<�D��V��+�y�O}�y�:nЁ'sL`��ú1r�c}�E��3$&�ꐬ��4����MM��NYO����8KC�I�9��N��5����_N6$bW�{���S�M�!Ò�����Cr&L��C�ܕ��>�>�M����Q�u�a%��@0] ��#�����ۃ�9�@D*��?��*�KC�]� �kG��/�Kl4V�|ה8���%��+��y��ŔG*��$����,_3��A(g�ܯRfHC<LD�7��{��{�-M�ӛo�6u�>5�';���٢���ߠK�57XN�X���u�ty/�~m�;
�^�Ѫ��؎8��`l��tn�T��E9�(G1��f>�Nw�-}%m���b߇���y������fm{�+��o,���T��ՠ�HY�VpY���D�����Ym}U���v��ڥ'.��z�[ᧁ���/f	EB]��oN'�'+�W����/����g�b��Uv}�������Qp0�<�����P)��jLٝw�����g�A�3O�R�i=��n/�%9'P;�XyҰg��=����\d=pfx�=���0D//�R���fF�[Cm�I�!��ʰ���0���w#d/SM�¤Y�nIia')iч�q�Cp:�`�k�1$�Q�`�@���'1���l���=��ˬEA��Îr8�K3�d��9�lD���@+��@I�k�;�'�a��♔���Vm:�ˉ?�i�ċg[t��e<�盯9���1�м�,S�y?��I1����6�ƣ����c1@�Ur���8�?�ll�;	������ZXKL�x4J�p�I_c��t�������g�?.��Om	'�}t�%X����������[�۰����ɴ�@�'^ŭ�׻ Z8�����I�E��}X��-��8�`w��=#�W��o��m"���$�� 9���i�������]� ?˃Y�~6̳uN�Z�qz��J�>�E���ZyH����J�[�t��ՖM����@L�9��U�֙��+�:�? ���N�[�7��y�
�&|F�������:�Qn�����q���D<��\Q�R�7m�E��o:ߗwۀ�v��#�E .qY�Pć�����E1)׶e��fr+���S������F`�j�l󹷀��1c!i�۱C�2&t� SP�m�Ŗ�Z�	��5-��:u:��0�!2^���.�"���e$lQ.b9K�F8��#��m���L'�)�ǀ��C���oFeA��.��s��t�_@�Ds�m��Ek�T��y�P(ȝ}����w�-$�Ś�]�D{}n�thF�eq�~��3D#K�
�ϼ\
HQ����)�"ֳ%)���\�����?���^�_7�����o���Y�
8b!K�Z��:`�[C��wpn��|5f�$�@��*Ax�	,P��D7!E����#�=�Z�eQe��i$�ڃ���n|C�	D??�Hx�T-��$���D�<<�P�y�INة�U8����aJ�5@f�[q����q|�Ԭd	��))@�9��A&Ht�����S��U��T�~���Ӑ˶���X��x��z��J:�ߘ��^]��Y]�DvD�la�SZV0�.ǲK��Yw���ٙ+Gt��%��>���F�G�!6�W�[j4=o�4�����4*(+��?0�M��R�M���˜�n׾�#1²[pl�sYr�>�,�܏���*d�KN5S愡0����r���I/[����r�vO��K̅c|i�L;�	<��}�t��">w�U��_y�z}�>�;@�񋘬��Ǹ�/����c��1�X���]�u�G��&Ƚ}��m����I���'a�I��$��x;*��~����z8�Ւ�k���Ŀ9ZR���N��Q��cX3��{�J= س��W�m��C-��'�����gu�W������7B}�OYXb��Fo=�Q$�_
����K���;U�ˬ�{�"=��I���H3�,x]�N͒�i��V�A��'G^�f+��EOJ�7a2�$V���ޤV�ẕ�ϵbJ�:�v����v�r�ኪ�ؑ=�@����Z��8�7��|�3w�&ďCrr�l����������Ja�_5*|����ܬ��P�n�Z~���Iw���?;��� �s�/��5��Tx��{������`���M�E������Z4멇uq����1�R�)��V�����e��0^�Nb�/����=PG����y���'{2�E'�Ț��Î�>�+�˖}<ΖQ�z������_ҁ����[/�&�_�r��Dc��"
�>��'�JS�7�Um:�~��ž'��X��ds�%�х��E�2��*��~��4�!�/˰�A�`�o�><p�0�v�64����k��5�0���Ф����" x�Q��I>��� ����>����OCE��F*=O��?��Gٌ]F�u��A�H�\�9ޚN���r'����UR�x��m��:��^�A��<鿫}��%��R�R� �"AF��N9k{ƍu��4#�RE�a��>�P4���6Y�&Q���Rm4�N	�v|��i�Uw{�Z�;�ܽ�K�(��/Ԉ�J��d^��l���B��4$q�����}�x>'$ev�Y�[b���ۓ�|�<�����p��0@��B�OG����[���:E�ܨC�\��
��1��֤�����%�'��ߊp>4�����V��6$z���¨�O���������2(�v��=hΓL�����&�b�؋# V�\A* ��V���?���˩�Gc0����Z���y��jǈ��Xi�-�K��`3��iJ��G_��q�{ƒ7�ɂ����}��/�,|x��!�Q}�U��<d��D+8��5��|�I�e�~��[m���,XtA��~����0!y��k6W~�E��Q�M��?j. ��i��b|콬r���Q�s�D�ğ���� �֏�C��+Աe�Bo^��I��;(�Z����0�IQ-}��H��Ȕ��6��`Z�w%����x7�E@ȓ��n������ox)��|X�&v�(��Q�4Օc�N�f��M(�zm9�wwʔ�Svu�\�D���[k�[t����R{�D3Ea���H�,/m����0z�YbH�%�vU�x�n�i�8���X��C����C�aU\F���(Pi�6Dߠ��Tp*���g˟3�*
�����N�9U��J�L���]���_�^���iZXU¿���}<źp$g���ѠM(תٟ����[��a�Z�q��"����M�@j��>����툌y��m(f&M�1F"�n��P����U�!�1�����`��q���*��3��H������C���j�ɪy@�@��1��f-nw��`�c�Kcʾ��vI�&^��ϟ ��o' tW޴�������W�8W+�u���$�>w���REN0�+Gk��|^�r]#@�3Ջ�5�6�r{��u'_lc�� 
^p�T�??�?�P�[�0,mV׳2��8�x?�����`� �d�ϰ5�$�%#�'�	��4�+a�==�`�"j�[+]A�	��^HT#3��v���Ck�n˄����#`]Y�v'������~���t�w E:�s�?�xK���M�����/���:���x�@�skh���Y�j�ղ��xR���X���|��C1��5lY?��Α?cx`��H
�|n`#(��KĴ7S�����xe`�0���~��xsS�TǠW�G��J�D��1���C^�� jUE�Lhى��W����ӱk�A��G<{@��j�	�KB���K�J-�d����	�XJ�P+bs`R�RQ�m���W (\���o	
�b�$�1�tu��*33U��W��n�~�п!�)���8�]�%��7����D��l����e�v��"1�7��k{�	_��a��	��c�g�ˈ������d�[�%�.m\T�����g���s�a���/�h���hN�ܧ�k?�E]���>�G	ڛ����Ѷ[���� �iSQU��9{~��%��pi�h�ᲟY��щ����SXL�t�Fs�m�� �K0�Q�6�&\�3���ŻX����c�w/�r��#g�ဟ�� qf~�Lw����Z1�����9F;q�����ֺ3h�����92�\347�t�Z��\���h���e"+��L67
�~&�|[���}�o�C�GQ���u(��5)��۞�Ò��]�G���8�q�:ь��,�E��O-�%=��B&h��Wd��C�{�V�?�`��"eB�HX���آn�Q��ݨ��ׅq��I���2ؿ��L)Y�?.�B�
��#�ee��-j7p���>���9nK1�̹+��MXD���E���L�i�T_4�Q�V���h�9�W`�_�r���'�Zc���8�G[2�Y^����V|c^��� �`8�ss^�E����.s����
#�!9Yg������_�EAr��4��o�
$�+�O�?I���'S	�������1
����!�4q�̋s��TU�w��d�k��)k�D�[rq�,��; {_���qQ��9c1<����02������r���$aTץh�U��;�Ɩ��NDJ��32���P�bC�8��%���l�<��%��ݽE���r���Ǽ�Q���7��E�=*�`�~$��1��)�-˔�a��S��q��`Uo�����<~�va!ʺ!��
(�2)Z �#R�m?��z�yg����ٜ�kwV�����	�NuR���9�_�w�Ԣ[�v�������M2x����Q��Л��.V�G�����Ak� OA�3d��K5d�i��B����Q�>���N7sv��U��eS����{Ϡ)��"����txo=y�qy��?�A�o������.h�i(%"=es_`��[Aw��Ap�u;��i�S~+	]k?L��k��)��� x��r'��)�D���_��Y�Z��1fA��0@2P�������f��C9��I�`��1տ����n���OӆkF���Y����p��ęv��WF�;b���&b5��Tk����h��	����~�_�|4� ��X��c�� Z��p؆4"��X�z�.c�	��/o��mx3�oϰy�ot��1��Ѽ<y�����` K8�?ވK;Ҳ�X���tg|o��ZZ|�X��%1�w?�d����rg��ƓC����ǒ�Q.���5VZ�W��~HT6��ԩ�70*�O`p<Z�6�/�wH7��Y����Q������f`���
��2�"}V��U�)�����<m�{0WK�%�1/w�y���s���`�2ӵnDɴm��dcg�ߵ)�E7RX���4h6�~�X ����?�-�Ff�b��T�z�8�G�K�!$nV��|��~ ���E�nF���I�����-����� 52�\�kp�������g�axe�wRAQ�:��v0�7�F�P���$'s�x�NP�t�^@a`�@�2�<6��S��l��`|��&�`�x�et���e ��휡84ˁ��e�M �X�����#�~�GY�oX��ᯱx,���aK���~���Al������6?Գwf��)��@�[e�Ԑ���n0�yx�8�?�V16���T���JM���Em��,,�Kh�+�0� I���S��z�S�ꌊ="gv(���|,�C���XB��L�y�K��c������i��ݰT�5�j�ur���o��R��}7%�4
7-����,zZ!%!�pJ�O�H*�y'Dc��l�z&��$�������Y$�,m�:'�`�?�r��������0=�P�8�}9�Z���K���!�2�~Ҙ��_�c	�3�� ��N�l�ʨ�&������llD��Eŏ@!�O��K�)�+��y�k)1�Ź�v�.�n���<S�R�p�'�q��+١q�O���?�:�~��z�\��H�)>dR���^��6e>�}�����vK��Y݊m���+��l�V��ce������3��BC�|�^^�)M�f�U�|�LY�:\ �\U;J�j?�����'���2Z.���K�!�L�0�{>��>	w��z<��L�GwK��r8q0t��^�$SH?��U*;|�t�A �%�㰬CoYw&��M�?����1߬��%�_�D??t�~P��d��C�.vfZ�w�Y��d����X*p0U�)-\���d3-�1�:||��Ng"���\ ��О�B:|�Mn��ɛfhM������A	���n����)�wV�)Z�u�b��q��q*�Y�u�*B�F�cW��8y���w�Y`brzb�2��fgnb�	�54�>��1n�n�i5󛿈v��T�1�h�j�ˌ	�*W(5�f�h;�5��ǵ���2\�ԼWo6lӆ��T�~:>Cq���އ����*�Wr�k���NÆ��,Jpw+�
�ah]Y�6�G����FZ�����ߥL%rT��M�� �bx�J���:��ٍ O�=�p�)5�Uk�n�b�˩��){�F.���'�kH�/ݓ���l{Èz8�����8��w.Z�R�So�o�j��08S��cۻ�x��s�:�;�*����B��.�C:!i�|8����*M��TU&�$hu���LQ(-���\8A������w~�3)kT��߰|���%cPn⛐t�5�����`JFZg�@yz�T$v��Y�Mۙ�9&U	�u�۵_[f�־G�F$F����^���X�[	Z���@|�F�IFS{�;����t����$T��z�]nTԹ���	-�)��<�M[�'���
�?QT-�#K��*������V��ej"�g� �\���Y5FD�lvlj:�m��A�m�5=^��ɪ�3;'(/�7B��*Mġ̰�DK�>�_�����P�(�FtnIi<��Q	]�����:�rd4��Y�~y7�'R��r�����Դr��H�֞�)�����Ao?��&��uC(�ZV��K��5�aT׹E���=7\G�z���`zr�*sY�m4���dY�ZN��6�&F]˲�ֵ! ?b�G�0�߭�\�D8��$���nמ(��u6�I��J">$
�!fҡ�9�v��V0^�đ��!������Z���!��0��KtL��=JI��a@�S2�./GM�c�_p��ώy�Cf�R/h`>���|�d��}`�hO�__!TPנx�y:��!'M�j�Ѵ��x�h޲N�gy�'�/��3�X��"P✐���C[DT����A��4ʬ�T���3��~��9{q`��)6V�Jܮ�(=3����|��=�� i%�O�bz������w.��:Y�ă���%NA��>�Wx���15�����\��b�h�~��**0 R`Z�}�n�%s��SR�P���$��\��ؽj;���p@hO,��k?�w�;�OԷ�E!S4tD�?��q���h���� �z�71�Y��ڋ�G�.��'�V��A�<q��������g�N��t�D�H�8H��w��bY#Z�ۼ��8�<u$��^]4��@�jEEk:� �0���fq�L�͋L�C�H���,���ڕr�;p�0XD����;qA�6:W4����QRĝ��g�SY80PPV��=��V�ū^������ �tBr�C�;�Qmݙ��62ϗV����C$Jdɪ}�_�.or�dj L���kF<��R/�:���g��bEO_t4�J�5�E���m�ˆ>��~�һ� s�ґ����Oc� =k���W�:�ш�`���4@�Y��l�����d��H�EU�D�&��Y?�������{!sƜ����2_{H4�j�~R'��+1�� ��.���P����qb�k�/��8m">.a�kRr07����Q"�{��D�g'�h;�V��{�N�$!���z��NK�qs��q�TI^���Pj�ZAEȝ>{flB����暔CY����G|�}.�M��@�ؙ;�E��~�8�>�	�(�!����/eR׺f�?*k������4�ق�
�����ǟ�� MB:�6��ƹ:�(A8O{��1����p�z}mlx�Ә����,˳7�I�R\�π��abl}��j�LѵmG�*&-r���J��#��4����jW�eػ�B�gq9�����7�wy�Eî'��B�`�*���)�~ �� ?��o.�6u���p�}�H�;F�I�$�ģ�d�(v0��?Be;W�¼�H���O��7v.<��_=PA��"�턖]�1�!�ĺF���/�p��u���y���5 ��n�����ؠ��y�df�;+�����~(����8o�h���n0��z"���w�����Ě��A���7�܎b�JGH%���lľ$c\B�,!������=�(��c�uk�à%�p��+}'����n	b#j7/jC[��N&s�� ��<ݠ9�ߔ%L N�y�_��Z9/�1�|,/z����S]����$�4�z��ʡ�@zK-��� M>h���R=O淇l�^,q����{�&��O��.kc������Da[��8���b��Ѐ�^���Y2� nB��*�CWi������,�<���{{��1�\HxDl�E���э�^̡���#AN���F�>�٪�D��xA��M�đ��u݈�Y��A�"��𗿮ۖ�H�Hp�����P�w�Ϥ��;D��\��$K�
�ςMӫ!Ԃ/���8[Ÿ=O����Æ��!�O�B.�H�ں��7qlv�������f����^-�`�0����LU�bPt �m���4��k>jf�'�d ��>� M�*�Ï�E�	�Qm{b�� /FFD����%��C����S���z8ĺe"<b�ɾ��CO!ܚ[A�딡�s���AZ��F>�#�/6  �-͝���:�D�p�x^���� W4}�;HS�kKnI�_X�w�2K{R1��{�aMV"�|��6�.�F�.�����l�f�?�B��Sqb'R�.3҆=��27�u�����
ݐa;
`�&�ͰZC��c+긖s3�B�-̃w�:������tϢn����򸭦`r�;�Kt�����%JS�?��v��1*�V�'�B���~M�vo{��Ù��BwC/�8L�嫝$1L�I��~Wsf���V�u)6�f3�~��<���%r(�����ߢ>Y�^��f3���@jK�i_:z��+;�Uc�_ؕ�����3�jm���==pB�����|G����X���y���ΰfp�0>��۸��8K��2D=Ѻ�K'fW ��q��C7�{a�{TQ������}��-���39����~U0H�f�ʫ=�2��	��Ssr���4`�|#oE���W#S����q�v���R,�nEM=��'r\�?��w"�_�/�ypȂ<�ŀ��!7S��O|j9S}①^Z/����o%[, ��(�=c���~h��/��쉡,�����|$z��D �x�B!�p�z���0/�N!���a2g�܌�̝o���Xr�L�cu�(�E�"���A���9���h�����$	Ԑ��Ä6����"��f��r�6-�d��%)��'Ƶ�<;b�<SY]oB!y�����s-�l���7��~5gх8E:d#iΞp?e���>W��=�Ֆ�u����J�*����)�Y�k��"��a��yF��f�%Xe~@b4:��lh��Ĩ���|<�]C��!}C"p-Cp\���G�whHa�ȓ�+9���||2�����Y�	����B
����5����5=���7y
��~�s�/���Ҍ\T*dFm�
B��
��~�U/�NY��I��z�����׼�u��Y�G�����n#ݗ�3�J�{[��,�7k���� �N����ɿ7�E@&[�w��;&����5�kԖy����.~��������k�`���Bḅ�<�	?jH�!,�>��# #+�OKI 7�ȕf06��^��).���/.�( �$B���o�f���<����Z8r�<��O�QPj_�aZ���6Rx[î6�(���S�MM��|�V�q�=�Mm��V�G���!_O��%�b�y�f���
���8��|�N�8
�g.H�K�U�ԺE�,qh�7~���9ؽ�4�Orv��q�-�)����;WhF��-����%@s���J}� �P��D3p?��X6�~�x�� 6�j �26��p0��<�E
�s���!<�cB��!i=��qJ,��ٚ���o�a�r]Dq>��Ƚ)ר缰k�ꁥ�؋�yC�Qm����'翐����3���Y�k�a�l���2,l�N�ѭ�.���"T$IB�׮e���b~�N�l�����#˩��:�������b��;�B��?t���A�a7b'_����&����p��q�%��y5�eiG���� �5m�x#S@�ZL�|6p��MDp�V�4�6�i���<:6�CQ����Pp ��7@7W+��q$R�N�sO�{|��"���"zR�]r���j3��"+��!���픗�[P���?�mw����O�+�fJ��Z�Θ~��擰�>�ӣyѲ)�o��0`��xf�Z��u�,�f�[[ҷ�#��e���X(j�T���ôYA�"���_���y�eЂ=Yd��fP�"-u��;2��^���`7a�9o��'Ow�U�]��Ku���5�So$�ؚ/ �a,M���j���j��%�|W��2�p�#��5 �-��,]TǷY�mR�hNPTn���E\n<�oB9o��)�j=��#�z���|�~���:��8
ƚ,��� �#��Ё����o,��=�_{�kp7���%kpЁ�4ב��6�`���8^ Nj<��Tb���}_n��!�>�L&`��b}$����;`�5�x�9��F-��B�E�Ƭ�B�����m�U8"��@S�3~d����M)d�� ���)�vH����E�T������j_�S��*
=����U3���(X�j�@��ە�9q����\�
���ǿHXb4�D��ᤷ�oU��H<0���������0�!u�M4�����OA6ء�ۡ����*�SAYY/I�怮e��O�c���%������%�'���xJԄ�V� ��	�L��$gyH����նY㵧<���}yHG}2�W�:PW����m��c5r�����#pe�"���z)��a��2�#J��/���	�^�ZP��\`xSjY�m�dCS�֪�L����E�1�0����Xl'ގ�!��6��R�r���~F]@�<mO��08-L]�T�>�+�t���×p�����8���;BL-�<Q�?v����J�p!��b� -��/9�tNE�O���dH�Hؚs��a���(-r�� ��k����`φ�K8�r! ��r�h����F�crL�����*C����q�S�E��/@Ŝ�A��ϟ\�$����c�\bz^2rr�R�*�-��[Z�="�x�B��+�� W�G�a5K�=�b�#Ew���������d:,~Lj�^i����o�(�b���=�n�Λ�@���,���%QE��|��<=Wo&\�c�0.[%��_ݟ�)�Or�oOd���J7�8t��
�E�n"(����S�(	��kͶ|i!g>0!��4����E2V�a{�ȵ�ZlS
v&�뮬л�������:�Y(�cXc�"xz>���?7~��Y�-�Yw6	�a���4�S����$1?����e�xHm�B������y����(�BВ���c����-J���L���H�K��]�/z�;#'�P��K"�t�yE��L ���\k����ޕ�R�nx���l[{c�.�U�;�-VW��t�+]�G�]��:�	�������@rS: R{�\ĳ�K`���Q�`L��M��"n1��|�o�ܕ�nw�6�I�lŀce�=�l�=��+f�I�)�M+�m� �U��L~y�<�o��|��?Q��w�8�2]<�,��$sB���Ӧ�%�g�-+�Eᰤ���k��AXX�ZD��\��ģa�W^T�����ˋ9ܻ�R�����=��FJ��8P��q��I��|:z��u�� �c���&]̄��Dҧɍ��8�ƹ�<P����ٙi���4KiJ{��~@�C� Mt�y��%�1�;�����N�J�l4��t�O�(�&�XC�(�hO3��=�	N$p"����s��p�������\$�a�Gr��9�҂'�y�o��<�I��� t�ƪ�9�n�3I��m3�Y�}�h��Ǳ��x}v�Lo��h-@�2gw�����)JH
w�U�jdr� e��ha��k��PK��BFh[4�WF�p�*�G᭛]��u-�쿽�1{��:W��EI2o�m��K3$Pu��;���(�p��3S��u�ު�Uۀ�ӓ*C譎�vf��r��l��
��k/	4��#>e�1��a:�xBh���C�6<�b.)&��瑛��.��Y�k���0����������x_�v0ٺYKŭg� BC5�\#m��ޕ�[a���o,\{��a"!�
xB�or��+�Z��u���іak�w/�n���*x��0�e�	|��LS�:��r���gJZ:q&M�����V�v^H	(�2����mތ u`~�>I�4g��@2����4���<5�ߎ�v��jҧS/����m�8��i��W�%�	����'�;��$��e��fK]��܁+R�lK�$��pL�VN�H�[�Z��$B@sp:ys>��ӵz](e#��z�_�Y_ yv�'7�a
�����F�!j#���=30�*�(t�3���1�@���ŦƇk���/�3��'�t	���o_����(ٓ���|,�8���Cl4��i�$�o�'I6&E���[���8�9��ZkO;ƪ)N>���0�>��d�����[�����0H���έ�w(�֭�z���Ź��%�$��j"xĭi�J0����U��T!1��X��G���d��K'$%�8��T�+�oO�[�?�}��i��P���$5u��ЏPv��5eZ�g��~�#d��Sǋ%Q����3m�cب�ݿ���E{�y�V>&���ք��8x��A4j�d�w;��%T�EBX�v���16�{�?�f`v4����X/R5rUCå��|?(���gP�B�-{�c��g��.\��C(�� DL�����˸�gsg��L~�&� P�������O^['��=�_R�{�'�����΃�$:��B^�Ӵ����m��G�F{=5����havǷԠ����\�V�d�����0�\m�}�<���RHY�qn��g�.�����(�}N<�îPo#�|����$7����t����^����o;��\G`PHҡ���B�|�����+ބ
���C\�����.R6�����8γd&-�흷�eC�ƚ8UH� �>�D��efHv�)	(MKeZgرŋ�Sp�v�?����W&��}�������.\��s�6#n��7���_�(��W�����5�Ozm��δvi����S1'ҜK�!B��㕴���*����gh�K��5 ���?�6<���y�?M�~4/�@����Z{��L��>'���k�u���Mq��13�H��܆S�tu[O��r�`�5lD$`l�s�����L�ʓJZW�F��4V�v�$R෋Z3ϑ�3q�����MN�5�k<�����C~|�ӵ�r���������b���|T4Z����ٝ��A�9>�}������X<�Clw��o����,�r����p�[췺��$982A�l\y��.7!���doX���G���bP�Ԍ����8��e"|w�@xn�[���ݻ�u:��}	�����
@o�0-)NL*۷4�^�/�'ep�MYJ�w8�'���=K
���"�ޯ6��2Ӱ_d�ʏ�M�@���3^����ⱓ"p#�%���
)�3[F����)>��K����l�W`7.ͱ���9K�D/��l}c�P�Y�'u���ix)Q�v4fA[��T��_�t��^��dV��x2�7ncS�����5��kC,�W�;<�<�;ϛ���,��e�������W��ҸT�3�P��Tz3�Oo ��1��P��t�}���o��əE�{�ob��)�.��$��O���C��j��(�ա?�"�'�-C��v�"�k�{C�}Y����'OoXl�m��@c���K%M_��l��U,��y�E7�ƃɧ�皼EM�+%7�E#��㕎jA��	�����&'J�r�1F��Ev�md$��K�m�-��^2��=�4����]m�WL7а:�f�q��"GNϛlX�q��͗ʲN�h��@�{��d�G�Qo'~!T�G.��7t�$��4*�쁹$)�3�	���xM�]��������w�T�Fa��8�RJ�׀�g639�kc��u�sP��e��2���ސ(OhJ�{\{(N���w��_��m->Y*gǆ�Ƅa���a�a/(!y���7���`��MS���1q��?�-!��p��E	��~�]�&&�
�ewL�w��$z�j7טq!ۇ���\|��<���]!Q�{�aK�苮�z6����,aA�-�[��#��1 �<���t�j��`����09o�Il�ynr����.��&����J����x�WN�V�^l�s��:o`��<�V�?g���o���o�iص��
�I,��A�>t�r�7π)Ȏ��t{i(V�XA�O��]=E%�[�(���=�3��#���I��?�a���5� ���8�g�%���~	w	��δ�3�⬧���M�\��.��Ǔ5�����|���^b�+Uk���Q���|2�Th{��XO�DXa,c��@Z?�r�Nzi����x�8���كV��yzri�)<���Q���C���oZZ��yF���Ű��-W٢ֱR���'@!UTO���I���T!	<��0&7�q$����
k��O�{.�Yo�/E�n���Y%)�Q�� '��k�I�u�{6P�p�u��:��S.�Uk^�Z�Ŀ:w�rV@�izܒ��2��S>�#����X�6�ȃ�;�Mf��}Z9P>m�A��J�lJL��'����Hn�T@����p~�[y7kh�ϚqS��uD�_�m��*�W�-�_���
�>.ܭ\鲄P�R;�K���-�������&�
~l`m�oB%�ś,�{�*���ʞ�J�%JDm�P���K���ȯ�kn\-���x0�h���-ND�@wH����|m"�yԒ� _���N�CS�܀������Cw��S����)�ǽ2�A�^^��ED�0�F��)G���Z���'�PWz|+]�c)��<f{9D��ח�3�����t�C�bC��)Z��/qK��9T�����خ����?݉Vњ[�7D���5��L8:���}d���P
Yy��%��E�|�2��= ��gء�.�h��IT:׮OVO�)ɇn/�� ��kV�9�E>Й�|��gǩ���H��P-BH��Np� F_g֮�v���z�W۠ݩ"�ݽ@פh�`�ԗ�)9�5!��OsX�����J1ˑL+�Ȉ�sS(8{��,~ܕ�r��G�[��<�2d�$��	Bgw����=2�Ѵ��-^��m�s�z_�T��ND��q�:)�b�O[�?�Ԩw��	:��ϡ�A��=�wc���e�#���' R�Q^RT)8M�휮���v�pq㞡��]W�+����efS�8H��Ulm��P̏�ׁw��.q}�*�A���ꢊQs"Ψ�K�=�lI�Ǎ�f���G�ḅ�����~-�q���\?��8|�)�YN���ﵠ�_9:D{Rs�ҟ�E�R*���8�nW������q��9*�T"nv��o3@�q�g	�]vaH���F���y������YOv=:��� �����|T_��h��`1б�Y��\B�r�E�x]�Ϟ%-��1�O�^ Y���7G/���j�u�[Fp'H��Wv�|c�q���_�~�KOp��Y`�ؒ�g囘��x��Ʉ��Sg�(g!�uPG�VS1D S�����΢��]ÆV�'ڮHP�G�����/�m������p.�ѽ���I@�O�[�Uf��#� ����q��N��c��؜)Y D?���A�i����
��E������\��M�q�D4��ڱK��z�;6ҁT�@�ߏ{�gf�*�1X��Ĝ��̪��<:���H�5�[ʠ��W�ޡ�4�%��������v��X��2@X��ze�B��ï���
��
7�/�����h����^����ߑ�vA8��5]9�RX��@��5$v D�;�B?��"��N��;�[�y�(GH��?p��4�J���W�
}�P-��xK"#�1
�8�b�+̯��<Y�"x�54���-e���V�x��_&R>[c���͉�5� ��L��T�u����wV���n��TϮ/x��U3��M����L75�5��0B�����Vg)�,j�N̽te	��yx�(��]r"
 hɢ�*��ڏ-W��i��@�Fb�ā�i�RQ���Ԗ:�va�$IL���z�~�p�֎�V᭢9��^��*SQu�Xj! �M�G�Wn�,����Φ�����.<j4���B��p3�*��ۯ�[)�e�F]:0��I�wϸ���*�n��1������b�ڜVЖ��>x�,b�}�g��?��s�A���\'vpU��=n�}���	RtS����XWRs�ݟ����ü�V<�j�U��&�l�[�`��}���d-��Μ+��������%���`��)p�ݱ�%�qc�N�	����\(s��2�Z���p^�19z��>��i�B��/E�Z��9
k6���d8�����B�e��S����ۆ�f�ZlJJ%��@N��Ϊ�P�i��}��6����? ���|������WU	q�$��.��C�ⲑ���>x¿��e3 �A�������me�7���Q�%�X�s_�N�����G\�W�����2>������#T���Ϻ �rϙ���DQ;s�!Ţ��ݭV�V7���u�n�F�;���X/>��vz�X��{�٫:}by��l�cw�2�lboZM�;�v]���=�W<��@2]�����E)�o�4�V�����і+;�=bh��
^�¢�B������~z�bNg�k�|�!�.��O���%��@��`�.�X�d\	j$}!鱱V* �#y�-�
׉�
��"3���mDs���0P�Tv�?cI��h���;1*�T3=�ϲ.���w���ӧ��d�8���|N̝_���orJ����ٳL	��|��Aʆ7��M׾{����ٟ�^k�X� �>��a_w�]����[p`��9���j����0�M^����dȱ�`�u�tCgk��5Ex$���{i�&�S!�{'	�K����
!��Yny�|�"{��֯�A��]H!od�CE�j�Ǝ�[y��
������d�����:pv+Pxw@�y0J�y�}v��C8����>{(@g�M����m���f;�f��Z��V�P�*�Ȇ�0�Έ)gЊ����/��Ox\�կ��J�{=ک8=�T��Q�xq�Ը*���`�n����;1�X��_�a/8��g�����]�-8s8�<�
�OD��?��j��.م��6'a]ӈ%���7Diy`'@� ��Gv�i.f��SM�L��W�%�pP�XW����χ/O�X������Oꫦ��n'w��G<����W��/���7�������wK���(4����#-(P�Qb
��҆c���U��?u°e�R�ׯ.����$�������@��5f/��Kӽ�q�� ~І�U�1�������t*��D�\�Q��N}�, ��'�I}�1������p'p����ld��u�1V[��F?���%��R�y9����$`��o�fsx͙[�AC�L����s�/AUx����ojRTQ��7!��'ț�]��kf���� �2/����N����e�7��m�혒I��߷~���f�) ~~�����T.QDsX1�͎� �}5ڧ�F,�:�ƍ't O�tt|Q���~DѲz�Ez���ro`�c�$	��x�Tb��	O<�֗%�y�e�`�"���nBj�kbP�e��M;C�{-���3��Qr�qHYuMt�ϥl�, �wg'��\��	zvQA3[A�a1�8{��'�*��p��d��B@���x4Q�:U/Qլ�w�,��	s�R�WM ��$��1H�T<��ܝ����z'i�t�"t�c~% �JV�ْNf�6�kנ�y� �|E�A+�Η�<s�ԕ����oc�L����g���b�ָ�&7��r4[�x��T���FQ�`p/�K!A-��P,�ƶ '��}��o��		����<W�ΌX��
S-%�ʐ�lt^���.Ab_��4�m[��T;5���=L��SN3‾T'6 %��3Ÿ�Z����9��X�{�[$�)�A�o�R��KPH��� ���~��o���@�������5n���>>/�X��c�j�߭S����c��_� ����Q��CD��2tg-�y�̍�1���	+�n4���}����┋��]S����!&R[ �(
�0�TJ��­���2��ݦ���7(��j�\y`B�)�Tu�f �	k!�`aǦ��N�?]��3`e��'t:��@�����n�Z9?�����Dc� -�¢��(+?9=q�R%��o����]\�^yǜJ�����Z���I�[���*+1ë��'�ᲺM~򿴭��[��V�b�`��\�o�,�Dt>r�Z�>���	;�'�jjBHWڻٽ�Z�v�6���$}Q��V�]<-�-T)�`�LH.q�E��>�����ٵp�㓍IEҽ*|��`[0�5��Ae�L�z:\��6���,4�ˣT�z˓_\atRƵW3Ϣ���1� ��Ց��N���B�rG��c�=��Gk3��V+��	o"t�5`r��ۚ����b6���j�E�'f�-����^f����{3�|�l`�Yj�5��(���(�l^����R�ǠcBJ6��\���vb��O\d�����;�=-��&X����N��M�=�Oe*M��u�p(�.�ŷ��;tS�´�*"j�SF��2qc48�JW(�)�Ҏ4Eʕ�����3��-�d�N��,�
o������g�8���ڲic7	���m�8BOMZ�d� A4ck�M�p�k�	��\���Y[bt'c˅�0�A߷����r0CC|O��3R���Ck�~�֑�C
F&�k�b�>;��l`T����/ɘ(Ѻ?IҌY5�&Tk���ü��w�g�EF�NmE}�$�JK�֙�v��)����+�ѡ�繗2����À���î���͂�:�3�q����V���]$zL��}I���6�:$n+'���x��.N���V��S�̗̉o ӪE]`�G7uvE!�����ݓ&����,�_��qW��ec�]�s�����Ȋq���[ݹ�nbC,�˯�7<�Sq}��1"����x���G��QP0�<�C�����v��cZO�'tMn)9�[���ˆF�>vAR�����D��XfSuk5r��B]?����7����CC�i�k4�:) )�5[�w�\nB�Y/��`;U���:0D`Ҹ3�� S'I�����E�?\q~���Rw=�F:Ȁ� ���`�Z��)�O�x�C^�4'�������-.O�6��y���H i�O��k/C�^�ZD+�.�hZb�Ng$#<�s0��T�{q� m�cq�w/�^�K4���ýXR�#u�4��c>��|�tc,�<�7>
�|4{
�=JE3�Q%�\��,�r>*�7Ë�9�@�*7#բI���Ѽ�g���n��n�$���?~��� j��A���wh�BI9��nc	%P5� @*>��Ku����<k�3[Gq��:o�0� -�L,E�����0�#](C�I�\��O��ȷe��$�DF}����h<%pQ
	o �'��c����3:�I�CF0r~iH}݁M����]v���\��DFo_�a���]�E)�C�1+�7��( a����b��6�L6����;s�I�i��ò�Zu��yH6����������'t ��ij�oDoz� L������E��`��hb��a$�4P	^�O0퓀z�66V�U�39�7���e�$v��'-E3���k��*�l^���R��DLH��[��j	���������h����?�^������u��k4~�e�\�Q�^��YLB;�\yƫ�����P@�ܱ��}�;��������gA���¹�b+��6ȍ�sPK�5`��m	��4�+I��1���)OPl�vg�hs�aB�s�dUG/L��xI�d��4<�B[�Uh(j�QŃ����m��  j=�}lq�:�Su�I񮼇	��^dDv�;���o�l+e�3������}�£^�F&�]L�ٜ��|��vr1�xJ�O�Ӊ��6��qҏ��m��ߐ�f���q��J��u�.-E���4Y鏆�̛�TL^,!�#M�<8��'ˎ��׫.�y��ޝ��ix�CU��,�X�cջ��:�M�[Ҁ����*�d`�/E�ߢ�օ�O�1�G2�Nf�{���6�G��!��yoɍ��B )I�����՜$�ƈ ������]�8F���F�'���6Ԯ�`i�o��Ot�#Z¬~��ֹBY����Q=| a�E �>z-k[��	��ם��2l+t"��le��������M���ܷq��������D�*��Ǒ�t�1�a�$�=J7�'��a�/��С�J�v��iN9��E�"�1�wC��̟rC���~���b~����ܽfK�:J'#0]��`�*`	�|Zv�E$��d�m3{��h�!����UC|Ncb��+��B��,�Ln���I�	4�7
���V�����_��,tT_������f��T�.���%��hl/he����V
L8�����oʒ:�ّ$�z��'k�U��9�4�4���G�{#9Ѻ#z����X��h/��,���D3�ّ��x��@^kز����S,�w��j��wl�~,��j[7}�L|kd佇��a��R]���g���\�_������N2��G!����Ab��ګ;!
eO!�ZF��~�)3{q;������<%�x~M��F��.Yn�IkbQ��n�ho*��~(�֫��a����ht�:��M�'��ZNWm�-4�����V~eX��?��P�_��-�{��Hey��\ �f�����N�����L��s-�����$��Fe�Cwߧ.��}ɷ��9����g��@2�0 �n�HHT!	�o�G���S��9h.��M��л�f����;��P����A�qT۾���[���g������'J�!�%�#DIWBد��x��N�8���u망l7�K-Ih�Q��B�N�@αٌ�n�>TH+��Y�F��8!BǴ��y3��O~��!ʣ�wXT�i���n�*�m�j��Hs_5��N��i�=g�|���`E�l�@rd�i�a�fkܴ.\X��l�2� 8n���huJ����n �֣�{�b��oa�-��	������m9ө�A�k���/��l»����Ǔ���\n�v3�6�"�Ѽ�#*9�4!˼%Xmݝ"~����0{���{�ł�e��B�4%Wܓ�)<9��g�C���S��r4a]�I*XS��fH��fRϏo���zZė��!նw��x(���Y���H8�1����U�ta�F%����ƢFq~X)�����g��I2��9:m��7l���bY��c9�����]�B�K��8"��e�:Rq���u�������ХQ�x���RХ'�O��{=�'������S�D��+ �ˏ��M&Ln��į��2?R�i�o�M����A(-��,��� �g<��խ�j	�%��8�P>wy��,>�]W�H������;>}�&ѹ���N�
���qd�[�./d��Sl�",�w	5.	$ߤ�s]'�u2iA%�gBV��3�ot��J4�� -�Kdm�#W�u�jN6�t��#U��J����wKT2 P&�C��t���Q���L|��S��L�j�<}�t�M�-����ou����;hsL8?owɜ<��$b���8�ɮbmW�̦W
r+h�4�,�%�m{ˮPG�0������`����T�IR��wS�i�,�ep���Q|��-�X��%vu��z��i`��Յ(���{U<C0�ŒmU�t�y�����'���L���H������c.P�$�R�&�^z��7�pJ��B��8,�4�l4�<�T�H�9J6�+�6�9�U|H3�O\h���u�I>k�÷YF�M��Y۾9v��o6�^��nu�7���{�X���[�뻈�>����qn����j��8�ܯ
RX�(Ƚ��+m��Ȣ� ����g�`�i�9�×��a��>?q���?���v��G����ɥ��w*�˒��跈ك���v�G_�����\��o�
q���;)i��&���B�����&/���זXD�~�Uh�"�*~�B���X����
��*b�㟧�t���{��J��]�b�Ë���e�e�h(��a3Pb"�MF�=t�?y��{y����:Z;�F����ߴ�mk!��/�l�5�&]��!��A\Lh������s��{�����^��*��6��u9�K��eb�f�|j��mb������m�� X���6	��Y���w��dR��IgĮH`�6S>�'	���r���z��7�G<�FK��<	BͫbgD�5���5���Dk�Q�7:`�.%�;Ju��O=�m�~��U�Q��X<�b��g�%i�)��; �����9-�a���*<n��4	���� �'��0g$�XE���Hi�yi��豹�v��
}m�W-�]�/���Q*:���*j*"}�b���,9%��:jH���ە��4fdN|L�>52���\� �I3X㴇h<��󰸎fL�X�t�'̿h��0W�1�lC;��C��qQ�'��W��{�(���B��k�9���0J&˶a׭�>ϐ������]��ǧ2
ٰ���bMB��� 7L�oE�>up��LW�t�d��s�Fܕ���@Ҡ�wc��������!�"�a2��i7�Ĉ)AC�}7��%a �@Px�֨����`���0���R�z�a!c긺���3��霆��8�\l�q�^��u۪	6�"����R#�Go�hn$�Wd�*�����;���S�䆘j~ԙz�>�&,�oZ^2�����DB��o�=&G��43#�b���J^���uv�W��F$=�Z�;�p�z���°��r}��د�b���,.��e�G��ȵeIYcn;����I�gG����Ď��E� ���⟀�v��\��
9��q����i����GY���aN�A���I���z�8-��8Igx�%0%����K�k��D#S��n�̧�;�N�����2E��}�	^�s~�#z���v�='~����_��K����tc�O�����qL�7�C3
� dJ�?���%#�(���:�`皂F(��ˌs�� E��`����{L�v
������E�=�#��'� �5���Az��l�N'[��G����cz�C'�@*���u4.��僇�����)2$#\��U��L&����E)�L�^_ѯ:��9�f��@��fW���Y�e@���^oDP�^�)x�S�c��g=y(sK��p�G�9����Jٞ�0�B�:�~�����h�����i[���3�N�D�W�=D��HCH���� ��c��D�XW��
�2��=��5�Tr<g�A����i�&ʃs�/l�5P�O�z����v��g���6�V#�~Ѱ﯀�eg��j���ˠ��
�*
�ݽLI�k#ɛj�H���t1��F������r{]d��\-klU�� �x�I��	y��t=P|7��U�;U��&����9��`Bv%y$��i|۬�,�+��[�6_g��>� ��W\f��ٷEv��,�����P���Y�Ɂ-x�t��B+e��$��7n�$3��,������"7ܒ��[Ca<��H���\����*ږ�������������m,Ր9}:� %h��P���^0ߢ,&�\-*^�5�m��4��U.mk�\Z��8!���&����WѦ�r��W jK�6'k>7���؉����h���,)�e�t�CJ�nD�DY&?����v���`�^!��"Q;��Bf=�@���=�z�WFk��y�1��^�-}>�*\��=NS՛2�s�s�qP��!�*�TrXM�/���{m��!��ӝf�,��(�#Ura��Y#[S�5�уjL�=~3��(y��gx'w�n�i���L�>��j[��ǻ�\kA��-��hv��6r�w7��Q
<jT{�j����G%�.�"�5=�y2~�{*(q�e/s�5?�w�������s_����E�}Oi�h�4֨��P�7��=��#��}��x���g�+0�{䊖��Q ��Imsl��y ��'\�y�S\����'�Cw��a��q�B��!��,`��tKv��LR"cqw��Y��Yh���4.)�c��Z.���*��}�&n��t�D�3�խ�R fFG���M�Oڛ�%#]7'"��O<4/�z��3S�7(R�;(����v��A8(��v�iv�MQ[�T�TY���s�UK��T�^|H0ı'�hcb�����B�h��G4�y���1�
��6����m:M%<?.�!E�'��%:��XE��V��o@`H
F(%*2�}�	�<tb.Ho�7[���Yp�O�2�^q:L/�;�uV��zs����YҗQ��A[���Խ"������J�YMv�p���B��&���Rlr���ݯ	�j�{ l�t��a�K�щ$�g(|���f-h�9&4�x����N���A�3�$�J�B��e$q.t1�,٣�>x�⛚I�Ҭ�(��Z�_��s��
���.j촤3{�����o[�O?�)'�t��f`��.0�$�T5U��]yN�S������L0}��I}�@v��㹩�ؖ%bT��3[��.�P8\�6:v��-)��|��)J�pE�^�Dğr�S����S<q%ET3��>rQ�9<�I�o��+�;q���L��TA�}��#�Cw��	r?X�>E�n1�*O�$�뺌�4Q~eWI�i�V���}M������I6�H�c1 a���gHB=�S-� ���]V�Q���� |{���|24����Y�/?J۳4���fv(���r���Axϝ��ε�:��%T�t{l�WC�%�z[N���X�i�I��51o�@��Đ_I$��L'�7~����{%�98�ug�(gCa�Z�LS���^�zzzl�{��<Z���X02io�k��#�Q�h\���m��(?��{��Y�C���H��I�$)]E���藢E{���J��I�L�DE�K���I�W��1� ~A��C�0��z�(¦q��e'����z�6�TpLC�5�|�j�d]�Ë��]�G^�jb쒑�ˆ��O�C���Cq�s%��*=�B�����G$�%��L�b���89U2yw��}�K�Z}�᳜�����Wc:����L�<���S19B79?��2ɬ�C��ڗKI|�9�gT'n$�� T�U�l[C7xQl��u_��	u"\�3+���d9G_�!X��$�&*�t��hA�Q;Nf6v�=���d�}5�ٖ�T�mPRj�E�AzfG�2��"U�F-���k�֢�+�2���u��L,��(	!���}q_�HV8	�W00IR\MgK����n�����J:�v��b2��.�\nX{"��ۼ~�%��\z��!h1�a��$�f�㒍ML����y��O}�׬��������w�k'9A���p���G=�oRC���qٶC��� �:��$��P����ClK�g/��r�2����xql5L��)\0|E�ܹ���:������ZpK��~Q�6�y'�*���%�uR������4��s��h��UZ�î�fF$��p5,��|�������T%�����ہ� ��^���Бl�!s%�5ɷ����.��yZE	ˍ��[T3�޿�"�^�Ҥ����IF"�����|hmF,��7-��xgI�a�M�#�{2���������ˡ�tp{��
v�?�I�"(~'���������+�8��W��[�Q���B_��7�*>�F�a�x���Ν<
&B�M���%0��8���<i���|�F�>e�v���~��˲��|�8+-9����L@��{�6��,7=���?N/�lЄ[�;��Z�l)�e9�М\��ٽ��~�Á����z��$`o"?����HO+Y=���9!���sEz>�ڮS�8�h�OC�W3
��,Ew��W_���"/�E�.�bM2��m"F�)�c]P��ei�:��e�*����M!c�k~��jU$�j�7�3PAk�$e�_�l9�^����F5�U{�̕��ii1�[�2t�F43�3�%�Ǭ�Y�HbS���P([?�zR�}���n�[@k,�7�ǣ~�81��LO�@� ݊�������Mԋ6��=�;�N�<�,�yFK����It�ru�#��l�����W◯�Yg�bK
��r�ڄZu��s��@�،� �����W�̦L_���Ӆ_ݡj�P�J.|��h
��_�h�1T��;��pN3�ᢠ7`���!ąjq���)N+8Lߗ`�KRD�]�������3c+�?�5�w��B}�U�EF<š��������u71�.P��-y8�+�G�0��!�g�*�Y��*]��.1����׵�F���%��LU΀/�sP�xw2�<26&Z�y�<���,|�e��&��ۛQ��*ņ�G}��+���[��1���ʫ[�xڅm\�솘�>�}?�7eI��a�@��'�٨���]I���:XГ�d�a/Ɉ�˻�(��on;aNQ�m?�O�T����.h������JR��~�j��$+z�{�[�vo��_�p���$$$a���]1(��Hu���ʬ�Y=���,�=����]P(Z��\r,U�-ɼ���-`Z���A�{�\��'�. ��o�U��ru�hK됎�x��U0����x��}���	N��n�����.��0�x�5d��cU����=�]���\�ZU�y�ބI�o�f��� �p@�� �ǙP~{]���ӊ�e�������`C�x{0Q��Y����fD���d3�Ii��U�v�ǌ)��]�8T�^�K�T���F�1w����H���i�+�ׅ��)kgO�dܘ[�8��y:����G����5h\�ad�f�pН�����)��p�M#��������^�ȫ%;�F��W��X�� �Jg���2��!�{���W&#/'����8�.]K
s�7�tJX=}�NU2�f�����ө��
�Y��:��&�$H���B�5�'ɐV���K,t��y�_�U������d���3��eE��>��2Zҽ�Vsz�Ε�(O��g �g噸u{|�=Xj���(p2k��Q�֛���N�:��l
W�,�k�l��b�R@��X���S�*/\���QЃ�o�H���rc�_�j�:7O�X�Puh�:��C�՟Ì��s���*��"�d.�8�W��;�Wh�NmA"t[�|{�ʸ���B1g�����i�Dƀ�@	�����8�q7�Ep*�vV`��K�]aO�2E��aR�rG�KƓ��S[� �8�˹�u(�$$Z�:��O�X�}��~Woχ?P�&e#�5���.�s%�,�����Q�3�T��	/��h	bot{[)��CTn�*5;������v�ykŊ Q�0�,��MoTa�3�f0C�#ǡR�n�@��ƍe�u��R�gx��������@���	��� #�,&�}��#�)(�tr�5�"�ҳ�_��Y�˔��Gj�v��i St�ʹb��@�zIT-�B�͟Q����^�m�վ�&�b�^��o3[�&D��5�)pOp��$�M��9���m�Vƥ!q v;X0�ѐ�I���4�T�pj�,Rt)u���cX����~0�w���d�KҴ`w�y=����O�\��'\�Gi�OFc}g�*���@_PU��v|�h�qЦ�<�O�P�}R��I�sC��ZAx��V���D�TQ�_���۲n �_L^ٚ(�e���0%�RpA_f�!xwG寇w#����#���Aߌ�r(aJP
�2��z��zj�ׇ�bp$�/q���аTl�[�I�2�mb�Gez��6����eʴS��Ҷ1zNFr��l��,�Q����<��=���2�����1�	V�B)P2�y�}��_,���#���▵|i���g��˹eA��슒�mߩ�ƟljP_9({�M�oex������ *ZQ~��k_ָ�pIgL��ekV3�0)�M�~�^�0�_DF"��A�B�zc��khJ��l��Խ��Ԕ��g}B;���G�؋��b�B���J���)�$�{	-������!#��8�l�xv��(`�L�yS%���u��d{��x���K]�J�!O �p�ѷD��aCJ���f�rt�^��X�jO9���c�t�e��o=2D�����W%Jn
}��J1��F�zvJ��t^}cg�T�,�m�%>2-y$�͍�!�'�EE.趎�ʧN��z�1	5��3J0P�/Ow�U<r/"R�_��o�X��>~�R��5�?�����0�$�!���	 XT��H�_�u��C�Oӫ�iR|y�GL׳���Q�K��lg7��"&:������\�(J0-"��$@X9�s�j����P��I���d�o>`g�C�M�$����ɻ��G( ��Ae��(�Xz�1&C_�`@���2[�&0 ضav�I@?�3�6Ά��zP;%6W���n�U.ѹ�yyЮ.4`L��4ͩ>Heȇ`� �8ǖ2��fAP�f:��A$��oQ@��'��5H"hA��U|���8��
o�����I�S��t^�� T.*��C���ŀ��*e�Ǒ<+'/o3���YW9Y��IJ,5y�dA������y�a�Y�Zc;��
|	���ԏӀ�����P�Q���MY�.=�Z��4å+M���@P�"��P_������D-	��7?�z�"�.�*��%akhl]SD#��A9W4�F��l��ڠ쯗Lg���g�*B�|�9f��������g�������uD�9�����$�?�}�Z�-儴ߛ��S���k�`z��X�%u�"��y�-��Wv>��O*�7FjU����L�x����Y�,$�<�D22WO�w��l]��#NՑo[4+�}�-���<��U94W<�9^��!r��ԣ#P36��ww��s�^ֺX*V5۩�琶Ķ��N*O,�1��^&:�KEB�ϗ�b�e u�΅�c�3~�W|�*�+���2�2PN=|��+t�?+�����B�!���,C����W=UӇ]��J'L���u$������H]1���78���8�KiH>\,hC�\=�*)8@�F��S���4��SY"F�RDy�:�o��!?���7�^R�����R��.���a& �~��j�`����k�@��COV�a�i�X�	^f�� 7W�n8!��1��G�x�AaLC�AI��h��)I*���9����rl���yd����,7�������=����
J��~�~+b��-IrNvM.�Ǘ�]] ����TGChK�I�
�0L���j=-�t�'�6�9[=�)9c3�{�
�/��~)^;$�J#j�����xb�gk�25��<RBMNW��ǡcg���/�&���������!��e���`���Fv�%� �#�+��Η7�G��׫zTA�!��{�|kl��5,�0I�>:>���l���A�w����u�� <�!fiF���D������M��`.ͼ�C�6�Vm�ʪ��?�W򧲝��>J�?�K��+�hA}b�M�u����%(�TQ6 A9
ٲk�.�N�cBm��x* ��0i�-�\A5�޽zeSy0|����@�b4��ll�#-��'U�ݪ�T�8�}�dU8�QE-rlӇA#�L�����I�)q�&]�*��'?|�e5.*-�%�Wss,+�EH.*yZ|��|"���\�9��]3!Oԩ/����m����t8j~�m��u<E�++��M��»��7�i3"<��s�۶�܁P	>��w+�v�TK]����R�;��W��C|Vx�._�m��<,�:�4�7�	e`yD���uFMQ���]@��c�5!��	�������kг���@���*Ь,��*���?ҥ�@�����a��Qք~���`d��μ �L��Ӫ��W�tn�0�"ޫ[�8Cއq�oB���퀶�b����s\T���ԇ��z�/�M�>Z�F�W�	}qHN5٩(�����L�4^�,�� gG��~s���{4[��h.����_�g ֭������x��5jy=��>~0D	��U�4�mQ%��&՚�V����^�ׇ;�P�֙�B��
��BJ2���f�c�}�(����XJ�eͅ���NΓ����ȓ��B&�gR*1eRZ�Ӓ��?f���V���KW��KO�2�%�|�&�;Y�m�8{��٩QpK���po��\�\�l2,\(?}Z�s@�y�����?^\�8�o!,��<�MF�I�;Q�he�/ʤ��ʮ�7��4ˇ '�+���a��O�:8 �.�C���E+ަ􍃒���n#��Dɀ����M��_��KVhJvT�x�q�W%�5��0�N��q�[3V�]m�IV�&��b�<�}����;d�ǒ����0
�*wx�x6���rEK�`��4�{P���%v��V.?3��|!�z��P"�����)�S� �_c���5��~"����;>�����#q�T=w�}xA����t"�T�s	4�)���t���.���hvq�yTL��@W��{G[ �dns�/��%=7M��Tٴ�6\`1
�[q��_ܛҕ"���ꦿ�ܖ�1�aWh4���N��Q��>%XOf-����'PÎ�̒���>	�N6X��]�Lδ�Y�)��vbI�wPU�^=��Z����h�\)i�9F��I�+4���k�h/�m/e,�~��&���b=j�A�M����?����Bd?��g�k%��*&��"|��(��v��V����P����o�H�-�[i�@Amwn�@oӄ���o۞��dlq���j����m�o�G`���Ѻ��Z���ɫ�)B��?>[�R�}���`�R�m2ְ�f����ss�tF4��I��Cp��c��o��/�&:>�hZp'4=��Ka`X����$�"31���d�����G���٪��D�ꩠ�+�m����n�c:����])%8�?�6��cx�):��<�� �wF�F_!:�,I�trQ4�:����p(�`\�;�vRV�[�~ҢN����3H�1�N=�hs��<H*�?b^h��0�g0QDz���=����U&�@)Ȝ��WJd<q@l)�����$�|����q\`�|o; 5���= <��b���B��K�Ж,{�f�YW��:wŘ��4��7X����0j��2%�����"��7�\PO^�/���c���U�Ա*z�-�@��,�q`�?/�̪ZK�4J��X�FצF�,�ܻG^��#�iS6k"�&�������m���\�&QG$�`Ŏ��;��ٷ)�1}�2�;U�l�
s<��!�ڞ�X(x�밓�~�lъ��:�6\���P0}~��^�L�l	���V�IK�[�B/b~�w�a��8�j�l��j-�r����y�|^՘��ae����C��i�\(����\x�]1�<s��#$�Yq{��J\f�m��S}I�0
{M��J�1Ә�y
��y9�zZ��8�N�0�p�D��t:��k�D~�x���}�Χ��20;�AR�k*IF�@6�*պ���&MD�N�"ǃF�Q7�P����&q�8����6pT?pG���Z�#�7g���������\C��~���r�C�ٓs--ॆJ��|ro�J���c�É��G�7��uk�bU �;%����6�}��B�5��X�	��L�h����U34�;�Ui>B	� ;��1��`8z��zT��_ё8�0�C�X#��,>�~[�}�Yk��ꀡ�$��a�$:� �F0�W/V�����G�6�x�������8�Ix��D�t��|4 �N�j�&T8G%�]��vǿ�3�k�񪍈�d�铊cve�F4B:\��?9`l")M�A���E}�����D8�C�Rm�zϋ�`lߖ�p����N�����S�a��nu��)Ae��EI��#'�X�K(��h�8�R�z�(C�>U�mO�v��"k�p���:O��H��L:��s r�=	9kb˗�=��u���t:��s3fY�`㉈d�\�ڼ�b.^E�IA��������l�	�*Z#s������q�����s}��B]ܭ*��aH<�'�Yq���"%і��M/�~2|��힆��}��	(>X�sG�Eö���`����v�5�����׃���/�%����<�A�-(��.����wg] ��
�r��E͆Q:�]���G�0N@�b��o������:0��`w�H�ϓ��R�U�?�j��g4!���VvbX�0\�3���P�������Ƌ#f4֚�[5�L�{�K#0�׍"�^Ĭy嚛Q�h�5�*Ŷc��|��yq@���o��m��Gg��'�ʮ|�e{=N�
4��ekfG���0�2�@ˇ_��ޡ������j���(`�VK�7�"��Y�R z.����U��G�
�d��yj�B�B�=,Y��L��\��[�A�\>��Gv]��If�e�����sL���q�N�pA�I<� v����+��V�ΠH��iR~�҆;�U�y���.���%���'��P�L.p���Q�}5��Hu�Dg%��t0>�F����T�p��p�|��j�eY\��o��!� >H�ofD���X�Sw���X��{~��6�d�ˤ�[F��F��y$�uP?5�*J���s»n�c��Wg�"�b4Z�؀�<�L������Ŀ�Swm�t�74��K$.?(�>��d/Q�r��q{�&v������~LPǷ-J�5�@���D=1���Bd����Ꚏ#ک����Y����4X����Hٶ�T_P���e;��p`T*�|���`yM�Y�l'.��ݑ��������~	��h�^�yj ¯^_X%7,�~'���.�^s��X�S��<�SƝ�۩xm1����B�u���)M�d���R{�qk��L����E��2҈��ŵ>SO��X��i�����&�~�E����`�����2��OBl�s��Z�����v|"lL�/ő��d@!�[w�F�n��ܲN�>��g��x1jA�;Ham��Wo|�}���F�ʠ��k�\���!�Q�]yޠ��ޯ�:dx���S�VH7�6��kE�;|�f��R�)ٶz������k�0!S�A�j2�f��ز��4���T:�)�S�<�rdJ�ժ>��j����0�o�hj1�Zo�����/طˡ:�z�V^ݟ� Es�6�lv8S���%�jGt�8�B�R��!���t.�:��rg>��	9Ӎ��	�(;Dj��ǎ�X[��2�4�3����LdJ��n�}Q�Z�^��l�/z���ּ�ONw	"�1��_p�Dۨ�D��ʘp� 8P.[��֜Pj=��:B�j����,93;�D)�ï`P�X�X�1��z^�2�?�������r���<H��/y~�BR��b��7����`���H���i04���S�"�_�+t��ۿ�\���_���Sl�w� l|Ql�=V��޽�8�g����c��f�7�heiJ�8�������?���@��Z:uipr�r���W^� ����MoF��DS��q��/i��OM��Kr��&n�K��m�Λ��t�I]\����N����ݎ�GM���Au�]����kb��!�p�%E\12�����'�v�bF�<���Yp���9�˖��?)OHxe5�{0�&Bw�Q��:Z��%6�|�d(���H�:E�`~k�&��-��>	�{du*5��;�����%��X]n`�1���D�����U��vc|խ�&��I:'.��ɠr�<�� �k���,�ٚ���$�U�g	�X$��Ԓ���g�w�c�Ȁ�[����G:�<��M�dK����÷��h~y�sA����
�l���T%�c��r�}
��.�����ow�F�9�4����{��.�� �h�ޑb�d��3������Dk��]qeb��M\<� ��"�0��%�j��kt� 8�3���Y��5�x�D�[�!)z�7�	2��B�6�{���[>������ce����������̸����WU�C�Wq�[���+v;���T�3��:1AEKg��۵a�RHoSD#�ͱ�.}�U��^ܽ�*dwM�6bb~��"""+���g�tO�R�@�.���rF���HT�?�2l��<���Id�:�o�:���Q��O�9V2A�	Bd���]1=R5閍U�>%x��ͽ��Qݠ��������$��R�zf����d߂3�J[[�]�j�Ub�CQە��JJ�7EMeգ�NcNVʝق�y���Q��'�0<�&��o$2���z�cڹ\=�`qDٵ��,�|F	�Ӭ������/�x
7�i�a��z�����7牯�0���x:+�6�^��rn�U�*D�˚�-�Z;%����]�g����aS��9��L�.ء�)˸{3Mdm�$�5�F�O;P��9=}�s�ΤP���)|��ɮ=b"��Eœ�b0����O4RX~�g���Ĕ�1��O��	�(�D�`�sSt)&p�*�1\78���-�3N���6�}�m�J������)O�������H�p��l=������$���9_���U]�@�K޹m��m�]�8�h֘�!�rגZ0b�8a�#��4�O�ې��K��9�n+`Aa�0ߠr����Q5�[!HK������B|�=��I%�dv��S���v��"}/�F�KL����ݍ7��TZK������Ea,o���z/]�N�jzC�{���y��D5HZ�Lx@� �p�s[���ϔ��[�g���^B�|�,��J��U\ %�uz(3b� o`��.VӁ����D]U���*S���^�w��b�g˩C}�9T���a몾��O5ݝG@�N���T�`˙.
l�M� �B�y>+D2M�u���-���BVu9�����4<X�07X<�]�;E�V6mh�Z5����ó��
%:I�O�4�`�6��gE}	�q�샡]�@�G:k�nw�\��j ��	�)m���;i��HH�H������|g-��ߌ�.�\���h�F�(�����1��ʐt���j����K�Z+�r���n 5oA:��v97˴.2B�Y�S1�Sӏg���bzA�fG�1��L�پj�?�G,�\^�p�4���o�?�"��;�A��d�4kl�9 ��S��Y;�+��s'���Pl�M4��L#jn�
����>d�7�G�>kJ�U'l�E`����R�t�QhB�Ѳ*f�����j�I��'��+�&�V���
\lA=бr��m�Z��t"�����Q�r�.q�`#�x�ݎ�н��P�|���Y@��bQ�7�?�d�4����sZ���IMjy���7��!G�H��4�H�&�V�����s|�v�����ö0�_�{SU��Ɛ$eMu޲����W2�_�;x��g��5�"9S2��]O#�OLT�"��U��ލ��yEj�$���G4�< �O;_��:�śbi��]�%;u+�0�ev�ݩ�.��~A��@�*����h�x@�����uY�ay�3�(	Y~��mu)⳷�d���L$���9��ɠkx0��<��尊(~��`��Պi������иt��n��_�"���NQ,�#�
82�w��}h�mnK^~�j�_J>���kj��14�Y�Q!N����&m�q+�_��b���7�{��^P^��0�T�!BТ�D{�I-���]F㷆)hfŝ�2�>�
5w�"�Z���Ic���m^�v�
�/z����+	���2���c:�fLp�5+X��f�)L����N$k(Ēj�B��F�N���5�u����&@ёL��=c4}�/��1�;*$/���X���_�Ilj�O��1��SC�ǋ�t��P��Byr��BD6<�Ш�o0n���#ʮ�h9B;��=Ti�^�Widz������X�P��*<��,���W��R���=_u��;��C��CbN��d�Z�_x���Ϧ��$E�u���Vh�]�<�=�v�r�ΟP�]�1�$Y� �6�(��� f�k,�������>���>���PaR����}&��M�3��O����6>��6�w�Կ��t.����=B�bx����l|dZu� M�A��[���6/TJ4�i���M�+���
�ʙq��-��k��ȏ��'㣸�ܪ�ʶ.�9�n4�
��d�R�LAL�XW�Mdб�S)��J>� ��4`�H��(R�b��a�%\��2&h�Wu��#��1�K[�4�B턪2��F���:��3��`�3�,�Nf���
���O��}o6��Y��j��A
`������t�A���yM�����8��{f���Ϲ�&���u.�7��xP1���e���n\g��{"1c\��So��8�t���Nbv� ��t���[�4j=�#���'� wK��x����ݴk(��ɘ�7h�)��U1�Ȼ�2+��>x?`FTI/��N$Ms���D�Y�i��+P�41���<F8�>�#.e�@��6`�0���ξ�ڋ��s�G!�R.F�=��N*ޢzH�oD���J��{�ؗ����TF,�?�/��F�8��֤����	 �2��b��*���L@�K~��h��H(�7�5�51�ke_��G�β���t3��1E������xB��<6�/iE\��0��x���e 9{���,v3D�K-�_	�HT�6�N���!e����g�%&p�:ܜ@�������g̝�!%��<-%�2{kb}�+'�y������ϫ}����E5<'���	�X~�`���W��e~��j�DFcK�Y���+���k@�%��5(�8v�����M���*(�Mt5ު�=�����4Y捃�p�P~��t=�o|��ӣk��9��@����ڗ)������S����W�o���s��MȨZ�Κ'D2����r[��ˍ�a� ���%�����T���ԜV3��RBP����#� D��V���fr�a��(��[���ː���w��$WkJ�/8]�ec��8�A�.�M�^�CJ�����7g �)BJ߳ �7�^���4��1mP��<t|�0U���u`�H�1f'l��^�"���3�'�arsoe���{�{��穈@a��D��l6j*����=j�y�E˻$���!k`��+�X-	oY��u�AxNx\D�ks6U�/j�/�p(}J�����ˇ5��SP͠��7(��L+�X�t[3ǈ��)�`A#�B�3_�9DJ��'����g� h�)иW��{��E'�`��`+>��}���w�H��;#�d^*�P�s���F�(����1�&J�}�~�yKN�<�?ǐ��wl+��V�HF�	��-��M|���5h\��ur5BV������� ��j�mE!��؀�����љA���C�t�H������J��g�5f����4�,c�]� �5�C�V]��WS;��:�f���P�!��/��1����Y8��R3�!�gg��w����ψ�����r��H�4���LM: IP~d��ߗ�K����D��I��[*�������7���+��6�I>g&C�bF_M��O]M�gƍa�at9f�S����x�k1���}Y�N�-���h44BNryF҅{��C��W��uw�L$�1\X��=#��:�����,�d�Β�F� s 6��z�О� 3�7(7��{��Z:!�ej�J�`��?�����>�<��2U��]��IE워
��oz�������������~U ���t[Eo�Bm��<@�F�b�%[��t�4�Q����e�n/.�\�y�C��V��6��_+��-]�a,6����.�>b�A�9}������U�L���֎�16�¥����z�B�%,�c<V]菎���#2 �$��-���w��"�ި�
Rv�7SL'��X�h�g�|���(��=�@�k�6{�F���?{X{D��l�=-���B�E��$Tb3�PKsm�;��߻O��qjP�w��XK��HB�r��N��o�^ߣL��1T�V7��aV�3���=FCn��mZ�}^�����v�0�s�OmK��Յn��w��<&���]�~����nn%�l��kXk� z���� ;��*F�\��m���tqG����N���&0�r�r��������|W_�X����a��1X�
�#�{�g��=��'c�?��ڈ�)��w����/�tq6�qؙ���h�g}��ێ=w��W�̰����<�,�oc���ّqx�Xx]*FK�y�S}z�z�F�Q�J��pa��n����T���`���/�0��L�_L@�1цtv���v�ق]VKw�q��7�m��Pt�^k���	z����+ޕ"E�e��w;�9m�`��Ҝ���60y~��̈́��P�T�^,��k�b�������BG��b�j��X2�8v����D����~�Ys��"�b�Eoc��H��TK�c܈��Z-4�� P�ϓu�R}�˸Y-�󒄰�SU,��&Ų�T�we��8��NϓE"6�5@q&���j�p����0X"�x+b��e�~�]'�Mci;#�@�G��"�8T	|�6��~ ��sn��{��sP��$���¿<��@�x &����QȦ�o�X��D��%�i�d*w�뫾fuEz�XQ?h5=�Z���IB�=�J2��,��F؝��A�Sp�{	����/��ھ�Z_{<t�MA��ޘ�居�V���ݛ)����������&�z�p��}I�9z�g_�Pj�����xX��Ň��!ik�h����+�؋�������yv��et�?��������j���&�I�<�)GI�\��BN�*!.8�[��-g��p����U�y�ӍE�x�����}��U�k���3Md��:�����*��2j w���-J��x���	�0���ҍ��=���՝�y"�Vz6�)@����:3	Ȼ�b5X�z�Ha�,+�Sj�F	�7��$�u@�=w�G��lo�3[p�t�A�sv1@���A�T �Ie_ynN��o��8�1��ڂj{i�F���m�.,��s�O٫��E�IR(Vق_��9���'���2~�C�6>�*+R#����򛎾���V��Pʓ_��J
�H3k��o�c!��ֈ3w�b�m���;l���v`SS�=�C����˺%��fY���!�3�O�ɞ�J7.�Һ��/[yvF��	l�p��buvFT�U�>��}�F ��V��M��Zh��`�C��s�K�lA�HoCu�G���%U1�+� �U3�M�P8p9�,�� 6���I|�]l��J�H<�'G�n�^?�5�9��zȶ��jUpjv}CR���Ou�ީ��S��J��9�'���P׸�_$��(�m����C>55ֽ�,� ��!s���m�l���R� ��Je�J �i,�p�K"��'t0�3r��!�.�O�~Mjd�P8*��i��
�f�63��JeU�[�Y����fm�GJ� ���Dx�x��W�.��z��k��k@`�h��B� �$�_龾�p!\���T-���j��Hr�b
���x���9�jcmc���o\�I�E�ă<W�:B���,�A�y�Q%9�3����[F�-Q�O��;�Ph�<��|E�?bB�z�v�~~)�"$E����J����,ħﶛE��}	*�Y�C/HNH��.�i���+��U?8J �-���ܼKv�˄��b�}�-��-Zi����z�=��O0���q�Fw\p�(au�%H~�&���5�|,�X���&�"���N�WR���e�o^7	wNB��1���ff����[,T���ɒN�~�+6�v۽���!����=@��:��.0��35n�c˅S2���x�tk�� p��I����p�ث��ģ.k���l����C�Qy�2Õ�Qk��;�ۣ�S�ͭ��'BA^�ę���]�
egi���Gc$8J�؃�C!�g�;CS���2�K��:��_l�%��mY#��,5�&����t�Z��h�6:�x�����T�h��Ř$�	.�R�q�%y�U=x�Uܻ�&L	Ƴ�y�����\�%��7���<9*�	/��D�`qLzLCW��F�=��&zI���iݴI�}hU�T�p�$�����zC3"^�"��]�&��W�U͕��4?X���kZG�V���q�T�#�h*hT��L.��4�W��LE/���t�O���$&a�����դ��q��W5�'ڧ]�1��Z���,�B�t8�EQ�������#��b��1���"dM�߅V��v2	���m,��9:v�.	_k�Y\!=c�Hd߾�[�R�3�Y4fm�b�l���P6�ߐ%�/�I���}ߑ���i.(,��_����;η'X%Ɓ|�O�RB�t���jR�sp'����*��-�;���u�j���J�I�mu,������c!�Z����R�b�Aߦ��/�p)I�m�#�JA�D���(�л�Z���X�l�E����I��H��2r�I���w�u�.�G�>A��t��'0^&�ƒ�a7��ScٚjT����mP�$�>�Oد��L7(,_�:Ȧ�K0CǞ�2쾲˖��APs~��%��;��s���F�q��^T��鐽����c!h4�I� ���8�m�J�R�pR\���>���hZ?XdN�]�~��8���&|e�z���(�ĉK6Ǎ=Rê�����(��'ˇ�#D��� ���A�S/����Q��|MU�p�������v��{b;;�G:��"���Z.0����g���ֲ��zf{�3?֗X=(4�}��5+,R�R1k���k�ona����$���W���˕�ޭ�����Z�"�^���R��P�N����BY��u��1F�E�s��?�oE�79�P���F; Ugv�-F��/�W�eK	����#�U� H\�^NYw�g��hjp;˄��]��x�/��I ��%g�%�@n��-�	��C��D�׆PԓM����1�S�1ۆ�W%���p�0�3�;d�D,)��5rD��	%��(5lc/֒���ޞ������K���b��kA�<�vK� <�jq�(��IQ����b�3ɴ�gR�M@��6�����X�Fٝ��t��
Q�d/N����=��,&/ģ�pE�rVc���u�r���A@�^���V����A:��P��W���1iU?<��0��p�ڍ��ԭ�EꝖ|e!���w��\�I����͡?���n6n�?	��A��t��u�ڰLl���͜5z"�I<hj4��1�1{p/(��P��XҀ[�\�w��t�;!�`<�8�f�C�
�C
���^��Nྡ����8�H��"T������w��i�+T�J���6P!���Й�M|D"�%���Y<�u�xR��>�?za���m�q���c�K�L"ٰ͹��Y��Oyysn�_����0�#��r��_2�X�����*��6�����AH�����}��|�d�f@��H犱g��o���⤓J(C�O.�s+r�j����6s�3=X|am�9�-$`����,A�+i|�|��G�M3qِ�饏�$�[�Z��|<��4��� o[}x�����G�ꡖ�=����ʒV�xp5q�B�L���^��h��4O~\UlѦi�l�@5L�{��{��h��&�|�;��f5�7	H��>Er�m
��L��r��c
)(����B����3imh��������aV�Q�Zwo��K���d<1�j����$-���B�����͊k�0*ĩU��95j	5� T7�B��쨏�����T{���'�Q���+Sͺ*�LJ*3x&��z��A�*-��ۺ�:��7i��tj��X���lkA���2�L|�0��"^"�b��s��c�,��p���>�
����4j��SQ���w5V;+ :�\����ԗґ֥v\�OBc'o��]�,�>��_ro03?��^8�k�Ӓ���s���P5k�K�#��ծ!m���z���SwN�}��#�����,c1�ԢI���W�RZ/w�wK��J!�_�����~�R~��$�4�I�V�X��Y(f���@�n����r8y>RŞ֌G}"`BG�Y�^)u���#w���x3���-�ۿ�]�"���b�f��#Ln��H�[�@��w��͕3^��o#�v�|����˴ s���r�_��>vu+�`R�%T��YRq�΢g��Q�d�t2�$+��@"���2�a�٪�������;���K*
�QZkjbF�Va�HH9�}z'A��� z����n�ǩcl�F��L�u"��y�x}&��2п�5K�4�R3�}��	�,>t40�EkBdNa��˧��S��i��FHz�
RlK��C��� <���I��R��������^D�Z�4�y�yB��	1���u��>z}��fS��W@�`U�Ц=�q>���P|�s�����/ �p&���Qӓ}V_��6�P㳍�&�a�֞`PF�����3��[�Cy�����O��.nSщ�M���	�>�Db	��OZ&�c&S���a���
gq��b>��x�)���O���O����l�5;���\BfBw�f��dg�ң�L�"X|�S7-�����h�	 Ld���Rrm���D0B��ê���En*��!hoq��R%�5k*7�8�/AV��[���a�yx��7a{�\oT�2�9�BL1�&�lEM;��1뚏��9K���y+aP�-QP=�2z�� U{�ٛ���#u�ј�d�q�y�Y�T��0*`0NX� سk;�_ڝk��i6�'���`��-Jd�K���@��N3��4žn'Y�e���_�2�X��/zj�GV���I�(��ۦB� Sd%�hzb!+���+�g�Z���0Ra�Դ��M$a�èKg����D�Վ�0�Un�^�?�W�\�	�O����܇��?��=�iEL���t�,�{���7]O����M	�% [�D���I�2]�g��g�=��v�� sc�a�-;rʰW�q�����5!rw�T��H��	=vC��aٟv��3�0�3�3S*ck����O���m1��W��|Sg���K�x��bw2�]]}P�s���o;;s�@���*Zs'6�VLCΌ=$��S@|�HåA8�Tͷ&��9��{�0L��.B��0���C���[��-�U%� aˁqI�&��[��I���ȡ���P/�_��2U���*�����S�R���D���O�]1�6�:rT3���APV5�s��ڈh
RLI�49hb� �`�K�M�1���5���&�,G��Y�-��R��	'�����]S�Gṗ�J��
0d~��*%�!�ÿ�����6�U��zeTH�<�7x��Ww��`��X��06c2�
���JXїֲ@~���(�pU���	����w�����7x���Q_a2�^��I�7C�cVge?x"9��TJ�I5�n�*�9YvFh  ;�e?Y�W�M�m�s�>��I[��8sAd�1៏z���M����H���F~�F�٥�[��l������!s�5�BV���^���N�&3�i�����ұ�[u���!����"�k�!�2�I��؈�j[s���m� ��7��pT~�0FhI�Ѡ�#��ro��A�[�������45@<�:n�(Dhd7kjө��~�?�t����I=������W{(�f��1�=&FP~$�����ƣ�/l^ԕI�k�/%������b�W�{S1�ٙ[R׏�so���[8�T_i��H��a#G�ti�k�:{eΉ�5�H�c]�I����y[Jz���QecמߕW�Y&�m|ؚ�C�	.�"�-~�nx� c��[��K�����Âo���W���@s�#�}:,p��;	���Z�{���Fۄ��xn�,k� �;o($(k�彿t�~��{XMv$Ѓ$rx�/ag��@QE�ܻ���V�#0���4�-��_��|3��P���ū"\��M���U'�S� �@-�'�<�l�D�����k����8e���G�����O�4�,6�'�q�;`®9wiV�-{���4 �>*ζ��
�$�tU���
�cz�"�ZrΗ���z>����:۪r�z���ӱg>�a��v��?>�Oo5-ϻՀ���7���
�yn!��Il�Ӧ�4�cA�M��\��/�v��F��p$��WE�(DԪ�Hx�t|��s�Y˵�*l>��9H�����k3����t���"�)�F7�[Ś�����7���tݯ�V�2�Rn(�^&[�覴�-�a�$��#)b�='.�<��
����a�E�):��^����\���|9�V��{dc~n�!& ��'׀���q�s����@���G4�?k����b���Ar���C�"��O6�B[6�<���l.r!�t/T�S�_w�k�큌�E�d뵫K�J'���YЛ�|bm��+Թ�&lEb�7nS����a����7H*?Y1�iGaw%����)-&�M5k��'�"�q��hp�]�����Ǯ�t��H�JK�;��8O�명�AA��*��i�G���AL�_ۮ���#��JmV��v�3�5>�t��B�]�`�#{鷺�3���c��s��W�4���g:���({�����q�PS���+�],���3�㛖�՟��?��Q�Ξ�ʷ�hF)@�	O|�>:`��?�@p�s�O��׸�'>�+�l
9�r�¢A��C=����ל C���`��W.����#i�B�h���%�k����FׅWݎ����~�K#&l�La�a�B^�^5ě'��P�`�s���ҵny���ֆ�TQv��pp���{��S+�����3^'�rQ2_`�-��r�Q	���uJ'�x����hb�*���u��c](���b�
���ɎI����FlE���+�ܥM��e����LV����)��-�s:��U�8(pYjs��&`Q@E����nGr!f X�"�@.����{�a�m3�m|������n���ajp4Z��njN&
�c���)�Au��@�O�(�s�]�i��~g
�M[���(yTi[��~��tN,�8��53u���sޱ����X������N������� ���/ ��Q��͝�ޤ�$7��x�d��yNL�`��x���/.b��a�)r��Y�l���Y5Z�U\}�0hY���y�cʽ�� /����,��Yܷ�;�s��Q�M�n��{�5I��s3����?ʺ�8k�*�"���1�x���!�jI-� ��� �z�녶-�-���|o�e�����w�J��{�4�����d
_|��W��<[��3�0s5}��w�8�Nx� mf�Y��wY����E+�U����TG���nį�"&�>��u���g{��:G� _�&�I9�N��\ew�aX$�$�X���y;�YiQ�Գ/o�R�M\9I�����׾�g(�O ��%������cM�Cx�-1Ý�����R?��C9��+�A��:!�/��-Y�`L��>�h�26�n�������>W��ogՎKI(1�c����OH�A��
�V��+/U�������7�ĩ3%�	�d�����Y������%;Qý������������M��*VKZi|���ɫ�j',�-�o��M��j�cJXliwq�1@�M�,�|<&����Uc�#$�߲��ї %�&��dP;��}�ɟ����Y���^CR�ɭ��	�ċ�O�x�<�ݯ�����a]G��_��Fh+#��vǒq�M��a=2)�x>�=k���I���+*AuEC��6�����3�t�=t,���4��c*x�l]�n�6S6���^/�q�������,�sJ�%b�B�RQ�3�Lȸibo[�6k]2(:V�ڏ-��;��m��M(>��5\-Y7�Wrw��K���Q۲��߄����w*��k� ���T�~-��Wx����5��DC�M+��Τ\ٓg5�]�7��еL��V��Pz��؛�cus<$	��G0kPoe`۱�4�đVp	�ְ՘B8}��7�/I}p����
�K|>mS�A�5��������);���n�f��2{��ټo4�r��-�{�J2��Ut����!]h/&���p�'�2$��641�z�ft�q�^��i��xkb's[5�S��u6��eaZ���q�&�$�<z�e#~/�� ���AX���O��1l���$�D��0�$QX,qU,p�P{��²��We]쑯]�s'�3�4��6`dz2�o(}+����>�)��	^��^�PC��ZO������&�������L˩���C����#ӖI�w�8�3�&U�#�B#�s;^�LG���dO-�i[����\��J&<�eB��&=�ὦ5��<��ՠ{�T���f{$T^���.�t��� ƾ�(M�b��n�+"x\X�	|V��/�%Ǩ���G��XL��)��3w ֱ2x1hiQ0�J_KG���[���/�RG�4�$�H��U q/7�/��\�M zd�ň��Aj�ꝅ�h�)���>� �}�����~�iz�mݘ��R�߮�U���pA)�8��zKtV���Ϟ&ci��ʳ��_ �ه�N��GJ�wc�c�W�Cn�x�3WZʲ%pCD2�G�^RL�{�]�:��a~b�v�����zOj��5�v`UxJS{@xLj-a���GE�`�kR���I��.���t�=�cj/y��-4p��~-�����C�xM��1�>e������.R��+��W�aƎC^����Q�W���^U�p���V�{cN��,�i^M��g�Wo��/�֡�'J:;x�z�������VSvG0���FN���7w����d��8��p�NqK=�N��1�B���UUp���-�뎻s�
��|#�j~�����Kxܒ���'���ɇ3V�bd��0��/z)����<A�	�������(�WC�gSS�[��'��R��Co��Q���/zl���N�$d�Y�Y�,�v;�R��%趟�H)���������sw3v�����VF,�������t�IF��[)rP%�#�}M�W��b���z�aU��VW�B�W-V�@L,�#h�u�W�J�:�c$ӄ�N��$�;z^v]լ/G!�Qg�ſ���GA�{no����c��&��O
O1��q�h�hF3o(�j�i� �lYo��:������|lb��W!#��NP��t���5�A��X�D����^"?��٬�s˩�cLN��[��a�����~U���ŭ�HMzH� ���8��`��r%b�yz*(ʀ*#T ��\�v=w�*�G�.�yB�*��T\����9;���N����,S�_�������)��l��Aԫ�i6��8 ��F�7I��V{�!(���o���Y�<�B��
l��V޾��u�D����}����wW4��M���I=Ĉ��l��T�#��߰^q�r�2zC��?eb.n���P ��%vC^�Bϙ�@�rZ3�#䬁�K}���&�xt�#gԒ\�hW1�;��}��]\5�L!��i��>�"5$�1�� �X
^�B�GfUG��!M��M�z©j��C��coTဦK&�����y���Z�/�>�{��o�C!�Ck��������� ���V9K����%Qh�`��&�/�x��ƀT�J��j �s�C�����d7�y,&�DW���r?����#ARn2�N*��1��5���|},2� :��$ O&3�S.De�������V&P��P|�m�J����uu�39��6s�[�Q�Ti�fK+�A��a�����X�s7�9�~�>�6���0������چ睷|�oa����J��^ml1h��VM��L;|��m*��Wc�>8*J����z5�0~Ƀ&i\}�58g���X�7��{q%�U�B�����S��t��%��A��Tީ���n-W}��#2`8R��3M�Ar�g��$*���0wY���6��M)�]/�s���׵�ʚ�bd�;�ygfj���q���*�aa����~r��A^6+�2�5q!,�N>�9ի� 9nɷcK�������繝ԅ��|�����BW�ii����wH1�����}=>*az�m4�N�Qi���Ъ.0#Mu��O7�ȵ(�甽e(i�Y.Z�d��d�{�|����]�{/{_XiY�m�H�f�ӘrA��p���ю>h��r��̖G�~!�щ�\�Ғm�w6�
�d@�Y�wm�|yY��홒q����F���u�Qu�n��g�<��b['��$���3���7!ͨ�Z��PKEͶm��Z�aR߻J�S�D�hK�� f0څ~��Wx@��� {����<�*T4-��~	��ͫ�]�9�XJ�*"j�I�����l����ӻi����f���<ͻ��+��x���D)�"�{I�ک%������\`�  �9`�H�&z��k�B��3^պ�H���x<��O���ބ����˨9�sgp���0��4���bPPc	:q&Rz��*�F��K)ҥx�{Stw�x1�O�߼�н#�������2q�������ψy�~�ȴ��rv�`ŝEޱ^3���@���3�=Y��ڒ�(8��F5?�R<f�tJ%�Oٚ�W����ƻ���_m�eMH���+��ӟ6i��>rP#8���4/�Ȁ�w,	m�>�r2� 4ņ܊�/M�0$��x�6 �q���51�sL�(��eR����AM>RM�a��x�S�0s�oE^X`�Tr���@�8���`�j�Q���% ����0ٍ��h�� 9{�6�n��^�P�/�rrI�ڗޢ��8U6v�.��۰��"�Ӌ1�� l�	�\G[�{$Y\z�d���#ϰ�����ғ]��'$#fJ4��B���ʬ`s�w����J�R�j�N�(qx��R;[����@V�)+�RE�?Qt��!HI|>���h��n����N�3����f�|0:%7nQ~��݄��<���3X��r6�U��~�pn�}�>Di��;l�=�Ǎ,�ؐ3:����^r �);��JJMhz��<P�lޓ��k0�fK&�}v�+�H=�[8�k<�y�ȇ�{�3��r��+�S��Y� �@��hZsk�m�?XOx���$%O7Z�u�O<��T��\�-ٟc�r�����u��a��������CD]XW5�	!-�7������C�ҎT�~�;�j���g? )��/;��H{@�|W�9���;���P�HW <&�Z:8���I��+M,gȕ��\H�����L�ӳ��d��P-�ybH!R��Ag�w�C�햡-zK5�~c��U鵛����/t��#L����zRN|�+[�,A�tEeq+g�0�s� ��;�Vw�6Hxa��f`N'UU�қ��:̵�y�G�Up����5S̾�P?�`	@�5��[f��,���U��B2&Y����<E�X@�mc����i�;S&�fI������.�E�L��K�������`g�k��g��Hk`Tu�e�}fo9�r�Á��ǫ$^�f��;,P;X�Sۙev��(t���v㚹ZL��u0�O��	:�@���4u���l�v����z��|�$|���bОd���V�i��h�d�2)��I*T�˒c����֡��2��rA@���$+�)�=�F�1L�5�CvH�d�1�8N+�_S��X�$T�=�aYc_d�1~�X�k�������҅�b��·�z�laV�M�o�[4�����9�/Ro�}mIJ��wf!��!'��k��sGQ��J�q��|i�1_��NŲ9z~%��^t�{��`L�ꆱ��-t���?��z�zy������+" ��m���3^���B��+1Z�|O� *d�HK�-?�_��yU�|����z�N�`�����`�"m��O��q��G}TFX�!#���B�u��Ө�k3w�yj�ٓ��ȶ-�X�,U��k�^!Q�)f0c��Q{�$]�����.��D������_<4ǿ�OE���}����v�y�v�! ����7<g���SLv<z�Z\��y�M�DQ�2^����lP�pª�$�b����OyT�F���::��$��}�ǖ�(���5 �/oe���"]��;dS�r{Aو���	͘v̝z��%i�E�]�ߠ��Gg����K5$&�|����}W&��c�:0U
_M�QbDQ�`���w�v>�ՂC�'�?�7}7u� ]�i�6���
|���g��ږ��h7�@�ۏ�	H�|�괩"0�?�[7�!��Q>��I���D2h�E���ՙ�k�2�| �і�ĥ�p����웵M��~��k8.>򛌟xSā�W���C�p��#}V-�K|6f~�z|X?v����-TFszm�Q��0�#��� ��nZً������kw�H��\P�/q�X�> �=#��~��e���^G뺜��m�fie�p`q���w~�5�$���B8�O�~OQ�j�;�>�n��a�H��gر¨������K�ҳD)���l�\�â��iWBR�3GÓ��R��B�|���,h�
�m_љN��(� _����	V��n� Ӌ<�J�T����|�Diȶ{_T�2U�N�o+] d�:#�_��)_���Tr��5��U6{�v�΄�w��	fl+����r�+���A!^K䄃�Ά�E�==�rue�"��
}[�ww^�*��+yk��!1,A�OGw��*	����3���ݭ5m����5.��M�G�
u�$ج7�TtS�H�D��T $���$���J}K>0�
<u0w��X�
�h�Gc��C� �����||΀;���C@'9B�x�8qR�J��2�ړ�[�My����叿��Taj��A�lp�)�	�:�1��+a���>�!f��,Eş_S�m���PL�|�>���${�"�nH�Y��L����nxOԡ��s��&��6E�+=͡��Ǔ(!�id�d�K���N^O�'�����VK�� �M��v����t$㡈�Y�<�$�Z�''Fk7�I�v��x?Ȱ���WU:woe �:�3YТjG�T��`n��fg咴������@��~�&��
td���4�&�fJ��%�:+q$/�UG����[�r��QQ*��:�s�a.g��jꕮ��h��K+�O��~���P�f��師���d�&^��	���2�D�&��{o�~����eD�8��J-\n[y�=F~ᴗ:��ޒ6M0�OP�d]%:&_���)֣/c*k�(�����Z%��S� `���:�G��3G��V�F D�L�:i�vY�c͑(�^@S�XO5���$����t��L��S^_��N�Ky��sz��T-ܽ��G�����|m���O�i�"�R��׍���gnm��l�]
=�Hxd	�eP�����O�f��i$t��oU\5��R�OfN�4�sQ"�SB����j�~��?G����Dކy/��/'uM�<��U~�q`jj�;�����!��+��w��|S�&�Vܾ�D#���ZA���x|��� �N��i��9��:��b\�Dv�[��eL,�����	h�ѮW)C�����p�����Zĳ�.PH֒�a��g�fK�:e�2\l=��v�1�P7@�G�vQ��}���#ݱ����r�i�kpQ4LL�}���m0�'���:g�w�j@��J��=����m\�#�d���CQ�g�+	%�3��&���s����	�<Q'hB
�{���d9
�і��o��oT�L����v���p+�����d���"�+�e��w��+&�-Ȣ�D4�!0���!����"|��O�����Ov&�au����8�AC�l���bw��B�̀���J ���ڬ��3��]��@���;1��j��CN�	.�GJ�`���u�c���r�����9@�S��`��GN��2~Q	J�7mΗ�o������1����w��24����������P�\����8�t���@�CM,��G�+�VMqtK#��� �9�Q58�_Zi���_FTW5j+�,KVP��1M\��X\KHy��<<Ϣ����u/=��'uZB����^PQ��kٱ7K����_�J0X��"g�;�?�����c=�F|�a�[�ɑ�x$axn{�-z�K�[G ���Ax�O�����|��N����K�ǈ�CE2��@�ÙƮ� E�u5��$�g�x;�	�%)@O��*f!Cz�n�����+���35;�v����9~6���k}7���ؕ���%5r��h��.�3dؤ9��=Ph:�s�آ�
|�]�t4���d����/�¼�V�B��WNgH%=p[�H��?��£��Cf��0���X�ؑ��s�e7.5��,��ŷ�!�>r���� ��$�� $k:!n�����K�_}�-+%�^��%X����B��e��%u�����,$��l��V�X�f��M��o+,�
�����5��P�m�J��^��8ot��W�(D�yFes��e��翬K!".&~lբz�8x�\{�$!���꣤cyDM�O[��*m��J�S�.�l�hw�\^�ا��>� 2�IS|��{��p?��'��v~Bu^� ��7��+.����>+=�L�2ޓ�6w�� �����,?��s2(��F��H��D@N����s�u�?W��F>G�L�Z	'Uش!�j���X��0#Ӄ�{���-PD�()!M*N̍�Y��	�^�/�C�kM�Ե�|�e[ܘ���6�v�ը�����&]��f��VZ�o0���	���Ҫ�/eA-�ָ�8�5 ��� 3��t���Y�C�����N�{�S%�s����[2��Jr'ۛm�jC�$����c|_����_Z�E4�"�Io�Nm巔=w��9��(�i�FcA$��=a�2���@�@Ny���4�m���c���&�_ʷ��\���!ж��bY� ���3h�x�����Tbv�2���pn��~UϢO�f��4���K��3g���h�@]�)o`�;wh̔��`A�˞�N�0��2W�j���2,�䗩4� �,Ww����[zy���n���2e杮���Ef�tk�+�v�S/�F����y
&������أ-+C./䪾�����K�]�׹&�J��ӜSS��\j g�Ùb�������<�݁\��ȷ,�1S���������c2|³�Z3Th,����Y� ^	I�w/
�In���4�`������xϱH��g���s7@��G��s,9!%�3P�r[*�8���w�:w�k�M��F(D����?�^ R�F��p�u�#�Ã�M��sk�����^ц�(m�G)㎻�v�(�'��RZs箕�ATz�
�m&��#��)O��_K�r��8��������%��V/w�N:�q�:�r3�I�@u:��t���?*�ז��S̾������(��
p���`Z�a�Ʒ�v#�s
�ӭ�ʱ�I�{Ψ����ưg�61�Yd�$u�Y�+^�ރKg]���P�Ѝw-%<9ۻR�:�=e������Ͽn��DQ�"h/�"T?ND]�a��2��K��\m��%0gv:9I�rw���Iy��=%�@� ��%do�C���H���wC����X��.>טRJ�Ua�o��Դ�A��I�1�xT��R��g0�3�����f*�P�k�4SsH/mC>\�V�F��to��g��EH��	�%�m�Tgz�8����>�3x��Oiه/y]���Y��翷e�nd]�S>���N�h��8��GlI�J�M�?U�X�I��t�a�F//I�)Ֆ�+���'à��|����eN�#����;{
����$MnM��fW̎�}��������h�#�_��j�	�+#ɼ8����wOw2�5u� !Ƈx	;��6�~���A�|p~�P��ݯ�	 �ѓ�cT���ݜNs�Cԍ�Z��n�.��@�l�[�7Lp%(';�@'vo"v�or�g~���b��>��7�*o�T�,͒U��?�B��t Ԑ��h"�+TT�r�W����SZ�����5⽽�K~N&���e�Xb1�RHo�M�i�����=��C���l;~��>�%ϓ���z�j�˭���I���	Q�b��4�r�,�A#z����$�-�u��1ۙ�K
����g�vPU��d�?�<ټ��f��7���$9�Kp�|�3���Z��s�O�3�t�,{̾�y_D�\6~�Q��j���-)�쁣A.�bg����P�v�n}��ݍ���o�*��/�FnLr��6E{g8ؘz��c�O�[��k���τ� �+~��W/=�6�����{�W���]�@��3��p/�L02��9 ���@��q�=�_S��2�;;�S�B�?3c�ș
.� ��^PY��	�^�t=q�K��nJV�O�
�O�����19�*��=�1���7���M
M��<p$�iQx-���kC��as���A����ON6(�j^����b�P)0�,$�[wh��~Kd�q�J�-�5����<��ߢ���zܰ�2y�VxwqZں�8AbҒ��d�<痳�2&Z�$��
k��uq��NZ8w-���4@��)��j�kʙ�-g�:ٵPtIs�d�g�\f�Ji�j�)X�:��z���J��G�^4��6���:N�K�(�KD�ꌼ��������9�����WC��f2ƙ�%7u��I*�җ	��2��R4i�ycҒ�]l%��rkʯ����՟+�_�b_�
��l��T�j���OE杹�1U>糽����ee��&��"X�������5	��Y<ζVb��H	�+�F��5�?��wpa���?Q=�)�	�������- �Y��S��:����[��yb�A%,)9bZ������ќ�/�/��ݨu����<H�I��VZ/(�*O��*�,Z+�^��㐢����d�j�Hx��Z���D��u�����n�Y��)A4�o��̑*��16�Y0�R?(K=1i����js&��s��gp�\I3S�%zx�w���=:����aJ)�aAઝO�ȸl�:�z6���q#y�j��t�s��"!X�����|�剴|��8$��� 4��;�\�Ԇ-��m+�Ҁ�m���m�A�]k��ȉ�b�/�u���L����C����zЯ`�eZ�t%� H�$���)aN6�G�4�1�����x�����ZT��%>yd�����k��l��f�������܈��5��s�����������º���`jq����JuQ&e�=��{ځ�[��(�J��O�-ԃ�F	ښ`�Vs���"5�6�J� ŻF����sd4����:�@�A�(6\��5s��k觥�i�n9��+�"��G��L�d�wW����6���%i�=�s�yǂl��r�� �c����r*��PSc��Q3�UK�Zh��+��v-�
��E�Y���cB��'1��#����5�0�;tڐ[G�����lm X�0���T<�oܷr�ZS�d}P����or��\�Jp�/5�t�f���Ћ�Z�F�|����"�����1ߔƲ2�R�N�M\BY�i� ��Z�����G:(�!�|�g�Sy���E72R��:U�����֋SwHnBM���h2~6�3T���p4�`�����57�e8�V{��3'����[n�Z2���a+dY,���(fK$%��N�8ܢ�3��aux��np��贈��;��������xE*(�EAma؄�Y،I����ztl��#3��L³l��XX&o�M�l��l���Z�:ue�����<u���C�C8��U��c<%iV3�c�D8��EX ����!�3�6UuQ�I��=�3�S/KIx	��9M�&�L��BG�4t iGz]�w5^1Ƒ���ˑ�@ђ�?t����;@��n�8��p%��@�%���J��EURd�NǺ�qD���i��3dΒ�\���:�m(ZC���D��BL!�G7��O0&l	�N��O�Ã׈�<J^�Z�
A��my_r�Uo��)E!�@6�W���g~�"���f��!�Ƽ�9���1�}�ŧ�Ӕ������"6�د��+ۊ%�|E������40Ч�zې�̪��7@���|�p�4ϙa��`f&S�6�]"�Ql�`�DAj�b�2q�j�%s�X�{�6����+�Ys���C�^c\�>}�yv����Oa���XŜ+��z+ZԈqMC^hV�A��J}��DIն�6۾�X�a_GeM�0�nѫ��6*��l/r�SV���oyD�f������
�KE)���
�`V�3V�/K{X1�\�i�S=��'G�v@\ĻF�Ix�L����>�?���P�)6ȤX���S�����Nє0{8�o�W��O�P8�w>��ݺ(�B���(��v Ԋh|Z�F��;(��1� /��w Q� 7�ݹ��>˜@�q�?P���N4HL�{�q#�pH����n'��4�Ԁ�C<6�{B����Z�����n^���H�ۇ���b��!�C! ��AyQ魗p-�����v���1τ��c4Wk0�����F�m�ӧ=�ش⺵s��T�m�[2X�a�JHe2�{�}�t@Z�)�mw�_,E��^Z��c��ġצD�K��ڪݤ+'�STd�t`;"I)2�jڅ3lkz'��$��4����F:%��Q��|'�iP���+�UUQ�:�� �;
�p�T<�"`d��t�Ǩ��\��H��Vh��gMzkJ
�ůD-0�P��EK���sw"�{Q�&Ϣ!Mޘ��51�3ה��7�C�Տ��Ȟ?�ſ�O��9�Vho�ܒ<o�#'˨E"���M��������4��`� ox.h�� �,��I������l@ ��L�\���GE����/�H���MS,j��.�Ψea9�p���W��h>*��Z��+$�@��+���]%F���ś�1xʰM��|�Nu'�%���� ���������)�5��%V�v]$�b(��*5v�\c L�D�þ!���y���'I�襵�Q@�U����Dsh.��i#^ȼi"��w8��o�e#p`�����u$�nou��|�g=�57��1��jǢ"W�X�3)�r�|b�r��X⪀x�Oq8X��^�g�VP[�{=w����"��
�vD��O?�P��n��SP�3��j8`�9"��;a�A�o⏶a���j�Eo�ep���	�H�3�����:��zTX��0��g�ƻ#���g�oK;��{j"=�ą��BSTԞd�
p�g>8��@���Q֋+��H����=u�j,%�J��T\c�/��ܭ�%����k��d��j��H�U.
�nb�jE��TnX�3��PD����G��N�Mq�� o��Y�$���)q�w�Zt�����r(��EK/ �>���͑[Ѯ��P8c�8��d�O���H�o��}��Up"L�J�ː�����^��Gɚ�@���m$.a>���!�@=�yNF��c��.��&�$ƃ��]�4MGmp�I�w]`���H��DG�À�F�y`�U؜��s_ ��B����I�P8��CƯ��)ˈ�� ���P�ިWh��oF�6��e,�L�CJ��"�2�H{7ޜi��c�Ɍ�5ˉnϿs7�rɕ�	�.56�R���fw'b�����N1�DM~R��X�j�ϗ0����5J%�V�Ϭ��Sx _�z/�A'���RJ��Jn�x?\��h��Ν85��c�A$��u�;�s&u��:O0�HW�o����>�?'�g��`J4$�2��kl���K����:�Y��)�뷸[���dP�(z�C4�����L�[�钟
ll���?�ބ�H��hV��_��m%�N�D�.4v�������H��+E�=�˃�[h���Y͹<��H��@����pMv�1`*��.IȘL{epzq��в?2R���<u����T�=ڳ�݊�d�E�é�Q,�]��m����7�(j��m���e�ͯR�c?LeD�����c�ݮa,�*��n�:v�%P��	�������غ���A�N�D��0�=� |@�r�4�6H?V��������!7+��W����D����&��cB���gijD���y�bcR��E�;��.=`]ꓡm��|F.�2c��
��	n'��o�
���?�O��>�.�̾f�����g�+���+�vÁ3���g;\�Z!ő�dN,��oy�Y����{��/�U�GM�`cA~S�>�}S������_O�уL�(��q�s����1p�����z� =T��Ê��,ŗ�+m����L����ٻ��f�	p	^|�&[�����k���g,��b��p���ƪa��ZAi�J��,x�Yߩpt'�1�mo�Hay3�865�L����:��WB|S�FT�[�{)Me������5�f��>��X  +�z�fRR�͙��Z��+W��Tq��5Ը_r2���XX i��®�������i�S�%�꫻��zp>}\0�����S�t�JQ~*9����O,<̍p%��l'����z��U"��]�~�ܡ�
0�þv+d!K�>������7�����F�It�,Ls6�};��X_�(S�x���t��'�?�d@���ХkF{�ԟ�E{_��	�T|��~CXD���8��4��=^ �Ɯ�g�\ ���L�]L�/޿A�����Fȑ:R�sN���I��	��\:KA����k�DV*�5ΞK���y�ɭ�@`�/��)нXt��U8rr�7t#c���	,�N�rf��f�*0�����&�`Aén��(
�4,�cN2�{8��_*��҆!@���Ģ�����~L���,P�
�W���m]N2����N���͈���d�H���4��+>0���$|���^J����׈�>���*������	����q�E�y;�M��p���[�������ȉ���~��<"�z~/���}��,b�b��Sp3�ceoΆ�X����F<�'2#]hfo�/?S��t[�i���b\mF�eIU�&q��N 7�z�8�ĊTq���Y�V�s3��S!�9A�J���C������f�c�˽�g;}4��PV	���]�07��"������V�x�x�<qc������{Er����=�\I�M?e'���Z ����	= bI��<TL��爔8���\�"D�FP ӣ��o��/�����m����(���*=��fl�k<�l��Ųy��]�:���Y�ىr�:�o���N�F��r�$=>���7�%
t��+��^%�w8�����H��x>���&?�iՆ�4:�fI�\�n�����=wC����"�� 0�x���VeO�zh��7����k��� /�pT��in�ѻ$EKp��-��������EV��ppq�}��O� lޫ�>4<���Iz�:gH��G�H�b���c�'���2X�*e�	�������l*�� $�l^��B+�g�WG��	�]5��^��;���
��܏���w�\�.\ܽ��uY��,K�l|aO����q��%E��&��z��_��]�)�e����>	�r���"�L�v����6)��-ѿ�S���ŀ;ΛQ��9����ӅF��O�u؊�481@]�ڸ��S���#�iKv��i��~f�.�pV{.�h0�0y�ѧ�����q���5}�ZS�Ч>)EE���ۆJݫ�
 �l���3㳖���k� ҞH�/�r|V���n2`Y��m�	5�N��4�r��=z6���4�`��p���R�m�Q �G]�+<�i��p�fȁ,f6,�Y�.J�5'�``���}���@�2V��j\Y�3��$>$�e�}v1�,��3Ex���jzp���4�G�#Zwۿ:�u�H�<1%�}u�wԼQ�I����>O�Wlq��?�#�W0{�AG%��$��!W3��q��2�cD]��J�Mi[�]���#��R~
L��8�����睿�9!Q� +��k���`�-�t"^���:+���yhÅ��5��t<J�\s���v�d���qS�
]�j��8<T]���	���*�K�ԣ�A}ӗ�h�a{O��$�.t�����(���:Q��s��|�m
�� )>�Lf ��`C�0�d�M5}��_�#�S�FD>�����o���cxT��1y-����:���|KC�1� �\��|��7��S��>}��ߦx�J�k��A8ϖt�������9��BE�8����q�AP�,"\����Xg7b��LU��3�Ԋ	�%�A�"úS%0��F��%��e����J6�T�R�w��(<��=S��#�����7�A7>��V�a��ϽTޱ�P�k+�5���%P�In��Pm9n^̐��ASS����KC��4�*;���;":^R��A�"���'�j�c���c�� ;V�r�ꔐ�K��a��~)�ˤ�'h�x"��]�+-�A���bK�ǆ�>�<|�g��`c8~�ݮ�t�@t������J��8BW�Y� ��@�8��E=X;��knEYi�Њ�#�,�W ��ҡ�>���d��uc��Q��d44Z^zR�	��y�j�7G����K�8���@(���3��\m�t���퐷g�\�+%+Ew�g�7��˄�̨Z���pz|���pnM��*������:x�»#Niv�׊�	�yR�S%�o�l*n�����ӳ�����ԮJc��Kk���z��؛ Noid�>܊ω���4��9��ǌ��^LB
yrɶR��`,�W^n����%�0�Z�'�ap٥���H3�Qf�2�ѓ�������~e-Ouuo�M-P�%;lT��d���)l]����l�t��Y�W�J5oU&K��(���
��r���Czs�'��	<D;��C�f�R��g��V�%t��_j��¼"R�3s���VgցCq��ĉ4�9I7zx]+b�8�.�#7T)�:���ޘ�6^C��hi�?�8�
:P�t~*�B{�$�2-�OU��m��I���Ի� � h��a�g�r�ml�hKy��qQ�����1�nx'L����N�<%f4�8�wϥ��@z`��ŐG����n$l����t]:�dc�l1��������B�q�GVr]��Ĳ��`PX�]+f�� ����|�9
���Zѓ���64I����$ܢ�MDju7�'V�j�[[������Z�D�	�bx ���R T��y)�6YP[�{�7.]:/4n�YC	9Z���8�4�B�f�t�+K��R�;���Y.���w���@|��|*K*G��2,��6�0��kc͠:H`�Lś7�6'hԧ2�Õ+�-ȕ���"ė��ͷ-�SM]�,T�L"�i�*��|	�v?�����l]�URU�y�r^Aӑ�N�x<�a�ta���v}XH�~���m�#%ܚ�N{�{�6'�+E7,��zࣉ�@��Ѵ���x�}.�2��h�h��
�Ȅ�����W̼�*KZ�������pBZ���$?:k�/� ���P���bw:�9��9���k��R�z�*��b��&�d� �>�(��f�f������Q�
��:�>s&���$�ꓶP�}�"��q�3��i���6���@޶<5'=��W��!�s�hO�MK�?�����c:�����)���$�Co2�Iޯ�O~�&h�eL�)yzV�f(֊��ҞV[�u������EF]��#�Zgi��P�2��"q�M4�G16z*�m"ʠ�3ep\0��Ķ�����L�}�6��	i��h�2��ШAm%�'��*��y��[>��P�Ցġ4nuV"M�}�6�X֝����8���Ui���.B�m.`3��#�s�ٮ@���s�(F�3��l�c"��2�=v����>�a�5����r}�N�emz4\�!i��8�&�C<Tq��=�L��Z����Xt�8�������=���'�%)"|+�}�"{k��eRX|~&���/5ftem����z�&o��U~�ur3����C��S���E<��靱s�c�,G�3J�۰�ik��������z`6���4vlT^��k #�� (�-�`��"J���F��z��20M�Vm�z������r�w���=�JM�s"1m�M9���94^����l]��vO*O}+;N�H������+&?b(?���"|%aBlOm�%1C�>Y^9[�~�I�%vud��m_��ޔ��N\ݼh�ReL�E:���R~c��"	z�p� �I������P�޵�*�ɢF��j���� �g"%hq\�t�����׭�N��1���r`V��J�L�~�.kː��IW�c��T+ȍ�Ҝ���+��6G8���$�P����x�gla�rq�g��qe+-�h���w�\SlX��l�P]��rpI|uk &R���_�2 ��q`�i=:З��`�t�b;R5��9�rI�C�%�W���iҸ	>�19o�b����y� �δŔo;��5߹.�+�d�0N�)�5SV ��L��t{$йU7&�r���'S�$�6x1�4��6�dc�����n� ����\��Y1Ʌ}�Z~T��`k�ME2j��6*פH/�i�����ٵ��w,>C� Df�7���\��Ѕ�%��{�J1/��uH"���������* (�0x���*������v��
	��f�fi�N�I�"VP��+�K?
��A������r(�*ψ]�D��]�@,2�����D�$EG��b��HH`�Q�n��S��b+��� �)�7��y�ꤥ'/�����ȏ"X���t�
@����E�}�ªǥخtiu_�>(��M�R��<�c36Ɂ��,,1'����m]��!ђ.�#6M����^J�P�� �	���U��YE�a�4`:���sw���*���L�ώ*zr�X�=�i��3���
-��x���D7ň9�Am����|�2�\o�E�gM�6eh�n�7�����R!-v�ǳ�}�a\�������t)����MV��@=l�$���;7��Ac%>����xe��֬��&����{7�+$WH�� (ilpB@��)��gdg9T$4;��V�u���#�r8�̋�-�8M��UXL����#��cC���af|�p�/Skq��T��G�ED���X��%	� l��f��������V~�_�W�j��g��K�%���C���*���
�HE<���oX��\P��'ܱ�,p蔍@��9����юQO�jvQ�:G��"UGY�� ��tu����=̴��kB�`_�o�a�;��k�	�wX���%Ò5���Gb����5�/t�������n�s��dkcI���G͈��c�T(y_|g��W���eZ�A��|�|��8��W��?�����	���6��||"B~���������ݙA|}��$aPT��P���ǹ�j�V��v3w����GW �G�Q$���_u��]�Y�����1Ϫ��=/��4 8��O�n���B�9ԫ�w�B��Y����KA�'�5lI���$��.@������z��j�~�^��cכC�30E�$�CE�	�˼�CPm��6p���k���* V5�A�+������M~6��
����܂�Hzu��<�#}"�����aY�����+B�7Ck���^c��d+ěi,��'{�k�I���<f�������gE:-��q��~�����y�1�q�Lw��X#�u9D"���_����~�9�jȌ�8���<���P���xS��AJ O_> �*%t_�k�L�֫	�,�b5r�J�ݮ�H|%��av�����o��@V��~"3B��G6����ۧg���+��`Q�@�%�/�@���-���
ǛRXA��~ZQ[ɬ�i+v1�\�7�:ﬦ�󴄌��fd(c�����ɒe)���y�u���@�dN��P��Myhy�Q���EMc�"�xX+?X:��\Z'�^0A8$x��F�f�Ʒ��C�͎�����$���,�;����N���A`R�'k�3�+��Nc��}مL]�SSpt�[d>��j��|��a�9e@�8��S%TLhS�կ�����c��@�\O�ta}�<˞K�s�;�
��V[�.>��U�b1D�<�`Ҙ�#�z�\6�x21GII�3g1<3�u�Y�	��AJq3�\�"j)��9n��ӣ��j�u?pT���%_Ӄ�'	N�qP)����6�SDN����%jN�9ڱ��u�q��/3o==]�@i��I���M�����D�x��F6k��_#�=����m�?��*��AVT.G�_u+!�����ka�`�pG�ׇ��ɄE{�zj�yք�D�����R	h��=����+�
H��/o��O"�ցu6�պ����L���P�}����(��f	ՒF����g=Qn=kS��}�^(@�6���8�j!'�d_Y�s|��\4]���'d��;��
ؘZ(i�E3�/Z��������vY��oo�>�g���D-c��.����x6	�G�y�1G0�e9�%�1�'�w9(���Z��:+2�	1e$�u()i�������w0���SL#hW���'<B��j�/��˧��Uz�_�S�^KV�(�h^��������M�պ�,�$	1�:�!���2���Q���t?�#]�a�T��pKmo�i�����[���@��&�.���H���z�����\_�i?�Y��'� *�w����"���|<,������!���c϶4�w��H�2cʴ4�Z�h��/��K�8��5�V(GE*��ck���#P����X�09haw��9��حw�����Un�8���l�k|�RQ��Q�o���1�m���ؾi_\�?�6%^�H�{��[��p�4b2�a��F�F���B&(k7��_]�F�m��jH�'ag�@������H�G)�-��#���i�s%[�U�)���t?��=qI�g���E��x�k�~֘��,h��WxU��8@�k���6��`O5ߑ�3W?�C���͸~X�b]�	{�%z*w0�d�m���}�G���IL�\�_ɚ��v�?E�6p��)�e�zf�N���\黛�Jjg�'�i{��H��� . �<sV�;�c�����^D	�G���Kps �\�f�o������.i/�1�#�E
�;�D�{�=��w�CU���_��/�2�(��N1�����D1��_Ҭ͘;\�=�\��՚\�RPn�u�p�r5Z]M���<�� �i���Uy�ٮ��s�b�d,�1�s�1����K��t!i�<w�g��<��F�'��@��PH=NT����z�.O�c���a��ͼ�$>[T�*�P�A����U���C"�����S�_�E�������yn��|NF
���~�}��P�<LOR9����E�emΑL�h|J�Գ&�~?,9�h�!���,�۴�L�:�
����LVيQ�b-��0I:A���Wk�%��`s�Y�-/�W��$*���Y>A�ӳx_��H�M��Wa=7���J 2��� ?'R��)|u���~�r@�c��u�~�#�"��<�~wʦm{���4��R�����ʑ;H��S�aeb���s���S�zQ=#^����Cxc�o�ƒ�����Y>�<e�46v�/�$���q<ut��qųz��D��ORN�#�1/�TtbڠdhK �_�<>���QLyIm������#?^k,��gw�Z�,���Sϩ��[��=��ide%��b��}�`��c��@�i�#ITK��CN���h�esԧg
	��p^�3L����� ��D���m-�TB>>�E��v�k��$	dk(a�꺣f��?���V���-fl0 7���X���Y.�u3��Ѭ>��v��-B�!�N�ݫ��M���1�"�����E��5E��y��󡐅)�#��G�F��.�x
�F����UU�ӄ�A�ݶZ���n9`��<���U���
-�*0F��p���$�3���u��lF%��@m<��\sG�]�/���E����v,�F��N(��P��x��pT�H�i��&�b����D�N�G�0��-�R�0wi��H��~r�*��c-gy�Qa@���`J��<�9�.���i�pb���2J&��"h[5u#�B��8M�QL�@�I�^j~'�(�s����^��)��ҶK��jv���7��츄��
�ɾG$�H��g����BϺ�?�ǷC����EB�%G ��I7a�R�y�l�^��$�a3?��3͗6Nx�\4h���p
[$�)�Ȯz �i]'D��gş�
T^o�h~J��ˆI��_Ī���fI-��
���O�'szR��"I}�暝N����T�{Ë���h4e1��������(X�����U���&�� ��,)q΃�t0��T�<3v�?�"�*��j��o���{����0x����^�������� �g/��vd餜Z@J�3��=ĝ)�r����ɞ��zt�}��a�\�E�s�H��m��-xY��[٫��4O!�n:�Bd	���p����ЕC�$]����[������yv�Ui��nWnoͿFj��oa��ӡ�Z�;o<0V�,�fuv��0؄�#9e�����j�di�W,�e�Af`��-�\%���`k�>���KC���ǥ܆G�¿����ͣ���ڹd��^:�6��Ȗ���g��7������teJ1����Y�hv����s�ܗ4j�����%��ORu6�ˡ�$�.����EB_���u�M\x8%!A�ݥ��V�B_�J��h��HX"</���'k#��A/^/���j�B�=��b!k���Qj,SϘ�^9���2Z�O��u�Kڤ"��r���	�f�ر$�b�z���wM�)p�d�y��5۟=��ȳ����)�������}k�=�"��ܘ2���-b��ĦA	P�ۚJ����P�� ���.X���<��v+=k�DH�S0c�9
CۍzI3u��<+�ʠB�I%6�#M+q�"?�T�h����UF�aI�fn+�B���w�@�(��;XY�D��nYϑ����X�`�J5�@�����1���|��K��af�)5/���k���b:�r�?�r�U�{�Ϩ�\b���Vg"4���!'\�?�]K�Tݔ���$�n|F��q��ݬ�Z�Հ��������B4 �〫�GX*���~cl�t�p����9�P���b�I�p��)��ezyU���;�P#�p�2x�)	i�ǣ#���W����/�G�90�P3��7�|!�ٹ�������y��'��d��ȋ���7A�%�}>b���{��\Δ���~�̼�qzޒ5Ա���W�}dċ��w���a��ʈS�K#v	Z���VxA�Vߏ�V�K벃v�D�r���*�V�l��\�C{0�[Ö�c�<�j��^čxR�!{�~���-�Z�q����r��b!Ė���x�zrw���q� ��(¨=����8B�T��t�ῧ��-�@�ړz��۬��n�?�"�:��w횥��?%|��	���t������ M�Š�W.v�^���*�s�0ڭ�߯ �������Ld4G} &����g�0s�0v"�Π���*�o��
��=��= ��Xs�c��$����󌶆���rW�u���,�8�f��������S�V�g�����?�N6%mY�9N�hi�`����.0��|�����ל)�]�fyh�H\{`��*D��*#���z�}nsK�'�:��蜫/q��:.V���jAy+�
T��ZM���������g�h�{�{�H�����Z��Ć�+��`c,�
S��R}D��4�I)�'.��ߜ��%&_IP������0��?� �4D0�����pX6�ނM�� z�>���?}?����b��m����M��rٛ3Ko?("����K�5�""V��*�&���r��(�F�&o��;�'�������ӛ1�Mo:���EU�/����)�z[��+�2i�8v���J"��J:�νý���ʰ��j�8��s5��v=ơ�7��kw+P��~���Kրsra�հI��W��~3�&���~)}�������ض\yo����B�.[��xes6|cq9<mK4��&Ѯ�c�d�\k)S�d��fn�u"��ގ���ѬQ@sti�m�O�10\+&ME-v�Ί��I��������zX���_\Ψ��{�Z�����'Po���J<��㪺��CV+m�|tp�F��t�B��t����!5��y�|�n��^qBg8��S�ƶ����5_F�|F�w��B9�߂sx��㇕�m�P2��Z���ҭST�,�h��ɯ'��)#��d�މ����;�o	v%?y^QMek�+�Hj,5��ظ��u��0�700xL(���D�8����7&'�j��Ǐ��n�@/5l`��,!��&	�Z���.b�fD�Fm�0["��y;�׀���Q4�*�R�K������K��aPY\9?;�U��hM(�Ϊ?�k��p7s(��^-�4#����>�/�7�'sfX.�DP�z��He�����i���(�!^�7�JuW![��?/8P(��?�o ��%��
|�~�q{t4��ғ��؀�<S�U�]]h��km�i�B^^ٙ�P��'�7,D�Nt.�.f�N/��;ҎG3���@qUjD��+Fˣ�`�o��UIa!����՝���M1��@4g�B({� 4�p\l��p#�^��D�6���� �d�^Q�q��,��!ED��G;�t�;eHzr�,��༂s����%BN=-�1".�	"�[�o��Y(H]�Ԡ/$��f˷1��.n�/���(��=���Qe�ZO</ic���}�/��Y�@nwQ.�� �f�)}y��>e���x �.�O�}0�B�'H8�ɹ	��,�q�py3��hއ���en��Q�����3�����e���k�3��z�̅5��L��Y_Bz �cqh'�k�T�I.2D<#��y~�Rq�DJ@!���{p��{xV��͍���Ԕl�m�Q�	��w}ͩ�V6w!���BG�z���Rq6�"���s�t�"�U����f������ܬ�"���뗒~�,&�<k�H�g�^�h�x� ����z��ϓH�hx}Rkc�,l�FΆ]7���(�~�͕hQ\N�M�:r���W�G����i��V���;
O���th�~8m���D��y�G2���,���?��k��
��u�=���+O���y� xt�*�*��+�1-92��F/V{oi��S�TҼ'�@�Z	��Q����n���Wl'T%�P.�����t] @�M��	�7�m��������yQs��L�9.���g�Lq ���	DH9���`�q�\�_n�Pd�mV���byR�#�Ssc��T�sh��2��_>U,�B1w�;���p��o�Z�h\�I�]�̵��׍i���f����+�p�+�ip�~�Ӟk#G9��2𝝀�_J~b �w�	��i<W�УĖ��"��$Ȓ�r���-�K�(O�ܙ��U��^�զ�9m�)k��.� P�rэ��;����f�B�CS##��SF��uK�9\��ӧ������*;�ܹ;�šMP�
Uo	B*�����I�8~�'����!�m&�[�yp�av}�lbG�⏹�]��W�]4E�ָ=�LP�-����bP�\�!<<C�b�* �tD�'^����o��[���XSޥew���R >��(��[�㧻�z
�Bt^��������E�(a�j_ %Rʊ�8yz~�:�e�s��|�#=_�,��EEVtt�ܠ@uD�w=����h˵�mt��_��6f���c��n�iVY;8�md��I6�qĜX�^�Z�q��c�'���!3�.�[+��n�H����k
��>r�2ZE��?�ច����R���`%��L�fqB���Xk�"�ʅ$hS���r�.OH��eQ0�:�`7�J�BA�cަ/qI��z<�d���|�#�kb���W��VnP��Xg8+�XS8����r��ع�w�9̤�+nJ4vt�U��#*G+�"�����.�@;��J>a�= V�<��^�ܴ2���9�s�$�J��L�/O�-������"G��@S ���8+`��}~w�.s�8d�Gv/�81�y����{r�#ŐdK���A�!�*���!~�Y���@�u�Kck�xǪ2�C*�e�z�4f�y���z��NC�H�jځv���m��]�io�zx(âô1�sT��S���k�&�S�u� �U�)�(�jjL$�y��cG-�;fk�N��,2n!���>��M�I�����h�7M:�ޖ,P³V��9�KC&�E��%/(� �,\��F�K+��1Ύђ�]���!w* `{�+�6.7o�k�d�#��l�$6�Jq��3�} �n�l�K3:��
��I>�,)��ޯ.IB�5�[�5�|�N^B����_��4��%{�8<{�8��^�ۂe���۟��d���?��Llհ�3��vxQŊ��럞Z�
���琢�ML���b��u�L;�'�kG�:e�jP
��v�<��ާ5iJ�i>&
ǣ�ƽ5?S�m�4�d�8���T�P�1�3#��Һ�"�"@1�,�ɵ<����zF�R��
����n�.;��L�BdYUry��|陠Y��j��&��	GP��)f�ߎ9��D���F��j++��i�����גJ�z"`�Xg���ŏ������H�\Q��f*�y]{����d�(%�d��\����Ey�	G��cg���&��Z���s����'�r�+u5��s�"��!GҴE�r-���6>��34�u�)p�W_ߍQ�|s!�sǑ��y6A|X,�_l����U�&����b�Lo��e��Q��}h�3Aj2�6f���!����l?����?<xAb_HT��e'&;�.�=�2ox�r�3�U��z���ш�ge��z|����7MF��i��D4�#jJ^0��6��~;��&G�rr4JE�+�@c��@"B�9,4pof�Q:�Í�?�m�t"]��<,�e��#=��R���x�5�%횒&ӵy��)eC���6e����E(�R%�
�P�n�xV5�EE\�~�(�W�����%Z�C4?�Y9�_�(��-]lI�_!��L�]�"ɗNd�I��Cz5C킄B\ܨ�������Q��3q�����ȸ�S�բ�:��� ����P8%��	������+4�?��c��*�#�3�.i�� �\ dv�٬Y0P�m���4/%�x2ٺYV%��̯O�����͔���m�Дf\2];���B��c��d�̳_��9nI�,BwQ�Ã� V��~p��@'L�h�K�*�5��qX5�k�!e���ϡ�nF����P��L>���h@a���P��7_�,$rЪ49z�6����b�	�9)O��6Q?R5���QwY���o�,��P?Z�.Y�BΩo���$&�\|?B�vB���������,����9�_c
�C_�# ��Y糇�А�'a>���I���)^B]F�����T��Iڶo.Cq�/Y�N���d ��އ2#�0,`����Ҕ�n�=�oڬ��l��vّӗ<������^�l#��$�E����vH�� ؜]��+1֖�S1�|�g���2�0><��"#5Y��{�Yƀm&(���׊�F|��Ƣ䲁�c=�y������9 +v�zQy�&?ן<z{"h)��_N�"�����4zI!�����3:�������w��!mЁ̣�)�xP�����i�Cv|%b/�A5�Ԑ��D<�gc��pG��@9�U4��5���x#+o��L�t�������z�>��^P;��3ٯ��!��|�5���|��ޫ�R�+�5�����1_���Ը�w��V?���e�>�٬�z6=x,V,�I,D��Q�g!�O���h-;DQ�����T��G&��`�j�����:A��>0� ���㓫�X�waz�A��S!�Lj6������*}}�V�V�m�Rá&YJ�X&^��MלP5��H�.���O��Rd�yNs��`C��"Ӆܣ�+��\vaHm������C�F�#�P������6r���.fH�R8	,�=��Y�����������R�5ۋ%X�02�2���t��z.�f8�O���zԼI�\��G���ed���F`��޽�cᛣ����C��������Gh�:+���\�Zky���H��R�E������[b�5_�q��|\��u���LUf~����P��b��I������J> *;�Ʊ˞^pN^ rS��E��}l��Y�)�)��.�墏���1�� M�(����use���9��e�@��+��7c�ʒ��K9:q��ۗY�b�����e�����[n )�N-��Un�0�����*��YDe5�V^\�e֛n�@�������n�O��G�{�vo�b�=Ӧ֜�.L��5���cD��.�@���k'�)�R�k�7J��v��+��$oΈ�U�,㋡xo �ʆ*��~��ڀMPI`��.�����`�h ���#o�����Խ/�d���4�&�<�
 c�ti˶U|Uq'1hJ ���t���#^08H�G=-���	V'�f��pC~�lP�
�曢�)T[:Y��Bg����B��
���mܡ�x�C>�B�n�/INExWoX�0�Z��6â�����qs�uzm��6���W5$H��@ԕ�����$X�ҧ݆�o�D'��e�W��2��a����F���D��Y�̩
H1��>�9=l��!�p͙��{ئ#=ϐ�,�eｿt�8_36��D$�.
QD�_�R И�e�_! ��F{�.��j�H���&@0��DZ1��U�,˦�㡳�����:#�&w��Z���uc�/Ƈ$����!���!=�<,~z:�d��^��P�5Mi�Q�?���'P2��ja!ãC
������&�R��χ�)�*ʙ���K�{�]V��\�[ˏ��=�Շ� xRi~� Y����n��Ø+�7 Z2H���^B�6���E%�����1�{��t���>@����!��6U����nS���X��c��v͔C�ŕ���́e&�0�w��"K�T������[c(ãER���yJ�?�}�7m1RZ�d��bV��D��H�\���J�h
�U�B�q��c%!�0�I� u�<��Dƙ���'c*��;�]�-�?EF�'S���dHפJʷ�	�>X�0���Dhs/|,�"0���R��MVWv�j��Ý�]����Ḑ���uhl�x�B���v�j�Đ����_x*H&-���!�T�e���u�vsa������_+���}��k�(WL�v�@�n��%�0���o�orR��<��Ԋ��E��xM�'<����`�V�%��vc�G_�'�m�T��ە�E��mK�3�R\�8�;�s˾�X�C��2��or�.[���?9	�K9Z��fs��!n�e���M��G���H��9P2��'u�L-=}�Y�<W� RR޽��jW�����|Is��+��4o��1��àK���yc��_��Z<�H�@���2$v䘷I3=''cQ]К���{�Ca�c\��rOv��`GT5ȚЌy�5˽��|b�k%RH�vE��?��d������[���l-R�H`��J���K%Z��R���;��n;*,C�ܜUI��z��^�X��L:1-�׍NT��/(^B=`SZ#f��I�F��n^e�gG�e��g<�Ji�u��A�{YI���Qu���� �!�q}ӱ~
'��9R���֤
�K�U�q<���Z��K� ���H}u���l mPP�s
.Mrm��h䬪l�qXx�C$�&��U�n��p���;�,+x_�MZ��|�����}-�J���\�Ǡ����J�\��~�\>�*����gH㛳獖��0���<�����4�����6x���� ��o���V�a:�݊���IC�u3)��4��`Z���>�g!gJ��r�-Z}l#�a�1�2����Ƃ�Ƴ��ey��nT�W}=��N��!e����D��Ⱊ��ކ�l��dާ&X�3�W��-�e��� ����4a�K�`?���O�Ѿ:d��!����Z��i�pG�)�.V(����x;4[D�?z}�N� T��-*aD��]���+g��6��3a	#jQ^,�]�t3{���1�<1�ѩ�Db:P)���;".�Y{B�y�ʀ5�x��"W�P+��A\��ѥ��
1`���$��ڲg6�y^#�P4����J��6� ������S2Ϟi� �L���t	�����47C�f�֐�/��m�bh
o�G�@� �h�7;t�O�Y"�=� ,^B��??��ڼ>���_�=��,�[݉z����/��?F7i^ �����]�+��y~������|�� ��(�SK�7u_��0���4����g��_�4�GQR�&hM����|�͐�hz��FYe��i��=���5ѓϰ��AQh���ht�hi��G�h��
�U��O69o[��su7�1f�h����ɇ0�E��]�O�w�R�:��+�|e�.Z>�XP�Dƹ?8vm�⤀����L��8S�Iߍ��t\ zb�.k�{�ǘ=��׎��G��&��[z�S��_�&�=�(�����Aj����XDsiv%w�n ˦���������N9��P���'��+�T���>�r+K�vC���i-�C��Yv��G�`Zݯ*�QLi�����,D��j�ϡ�SoOh��2n�kFS�U�~�AKMľ��e�Ŕ��ˬ�������uAI|�eq5�)�	�O^�_2hzPȩX��K�<�czS���.�+��`}��#h�ʣq���ʼ�v=(;af�kc)A	�*��q�6I�/g�3��� ���$�3e����ռYXaK�I�)
�j���&I��=�&��W���j��9Zё�λF�QL�F}����9��Y�#���ZcxbR7����g>��!�
������\q�m�u��L��.��9w��W����RA��2߉�>�������34	������3�ō�L��8�R�$��NPd|�)fO�ƺ(�ݣG%ʳ>��$�"e��lO�`�Z��~w�~��>�U���F3Z��1��e����' [��JC3�E�i4���kc�BrC/1v-��xOR��i�Uўii͓�ϟ�n�I#D�S&��+ǚ��Nm���	\;�Hb
�A���cgH�8M#�R W����N]�ln:����ɻMB���Ise��a>\l)S�b����S�wb��{���Z�Ȉ1c%�.G�`��緳Դ50�� �HɎ0������CTE8���K�
�!l#D~_����u���y�N|5���n�z��y�7�g�:W�`\LS�d3f��bٿ�1�C���5�CZ2���J�ϴL#%ey5���T�{���T��2�E�Za!&/���p�P��|�](����݀`�*�H�xb�8�Ɠ��$"�4}���X%:������� �|�'��\�4�FyHH�l|�0�����3f�`T@�Y�}{�ŴR�6 F��`��TX\FUf[`Ƭ�J2|�a
�Hĭh\av�6`}Ni}`R�D�������Fl�������Wi��m6�#�� �!(]&r(�S���0���Hv$-����B���/��[����H(^g�!��h�JG�����Ԋ�bjC{�e�:D頻4�f��7q8v�WJ���3��feQ ��WJ�p_X~z�/���*K'�]�螵��+��?` `¯��Wm�i;���¸�ãLЈCT-@�x����.R��W�����[��~"Ͱ����9���;`�;`:3��.zZ��ՅW�bE�ب}�r,�Ժ��Y]�/���l��3�&��LQ7��8����%�?Dr�.�l3L��uc��8Q(T�� M�m�g~���W��Dۘ��]B2�\�/��cs�^��v?�m��6��*a�cnYP��nr�MOH{]M0�6�<�z�ڽ��<vs䷔���ؓ�`�NqE}%-�Y0�s���Cr� &���!���I���~>o�^:�F�X,���Q*��RV���
%ß�ޤ��x�������6�Q�.�����t֋��V�֓(uw wճ��V�����6��3�)��/�ݭ�7TC�Č�vq2Đ��=���Q�zF.��7������"�K�y6����(�{�'k��Z�V�c�_��Y�\���s:��4ϟ�-Z���P��ƭ�q���Ø�h�/�^�����T�M�&fƮ(�A�����r�k��-�N���md$�[�L	[W^eBe�ڝ��%S���̆z�� �����hɒ���� C��h�����8>�u��z�f���|v;�*c�Qb��,sy�ݪ�&�}3Ox�����)��ZV嘒��츹�|��̯�iZ�w��c4f��i!�,���y'!x���xਨ�o��hB�R�/�c4�����[�ĵ#�P,��1��WA�IOo��c����ӈq�����r��V�w`�J��hLhz��[Z[
�s�Ӂ;�V���\��J'�Û1Ẓ>�"|���% VZ�1/#.&B�ɐ�^��X �nU�ˑ$
2\��q�n�d�4#`���7q�,_���F����C�*���L�I����&a!f�J���n}3����.B�X����ʛ]��0�&/����&؏��TQ���&:�+�R��H�1������A��J��{nTj5'iw �S�}j<�z'�@$oۢ�'k.&n��U�� :��Q!��3�n~�$�:��M��E�t����dpu��h9篽��9 K�9��kD��א���;-8|��SDf>�d����úKDQ{U�Hp�u�7�DU��(�Ok���#G�����>�m����+���B'���g�I��G5��`�]����.�?�	��Y�[G}9��W'M>o>�%C�`QXZ:�T�[S��(q��P��_[V���+e:��:8:�EO0�T9���e����PӽK���8ܤ��	��Dh.�a�p[L�h[�*2�ʽ�{�k�&�;� �����Y�h�1HE�LOL����Ҁ����< �!we�\��� �Y�K���X���H��W�v��9�lf=,��۬`UT��;­�2��;��;�:���8�u��}�
6|��M��ʹ�Tt< *���Y����C�}F���C2~�o�D^���aU8�V�~9��Hm����󋗍���������Ȏc��=�cV%&X���z�'d���d��G�}���n������C�<�ȵ.�тF<,cp�v{;���ZP�7��r�G����=w�˕Y�%E��*굛�^���`@���^@�Y��Ҋ�c�2@�1迷ڔ��6d��d�X�,Q��"��=Y���2���:2I�k��}T۴x7ኧM��hW@s�1pr��	���a�ۍY�����Y��sFY�.f�L�|� ����v{-���հI;���p��ﲮε2r*�D��W��5���0�+4_�r��a�"��o��^Q)p�=c��gA��ZW`�p�=��*/����)���v�R�
������o��N3�\ԒQ�ɧ
�������e�z��&�:���@�c[�$[�0��3�d��dz��(*�BYO��k��ʂ1+ e3�S��l0zu�%�ġ�R:$��2�X��Z�:cbz�@gݎ��ك�8O&AOl��S�}���n�(���D�C�.���!K���2���N���cO���9��z�u#�uW�s��BV�K>�F7��̠Ś��C�KC,�� ����U��!�lS�*x!��#�'�_<iYǛ�T��A̕M�������P�xC���-HF�'�u�$�ޘ�Sg�
~��,�u<t�As/ꗘ]��&"����/Kn�x��f�٠�H;��<>���F�? ��-vp��X�9�7��羉 �}�pphC�!�n�w�*VW��b�ͱ����=dθK�����A��K��
n5���Ji�M�J4��.v2:Z��{�,o�k�h����[<���́xX{�m�ɸx;q��o#�R�]��a�O�B��]W� �&*VY��`�@��gP8�	[�1����.)W 3Ӌ7.��m�i\Z@������;	HA��\s��C���=�����K&oN�KS���ve�h~e�MNv)6O��� "q�/�Y���o���?�l�FÍ�,�M EY�����y��"UDۨ
���K�5t ��R���h�y�-�޽m�4
��5��o��-Y}���Ƣ�D+�ɵ���X�і���>�0(�D�����󩗪�5��(CnZ�Rt�+A�X���tsv������+J��\Y0��)
�3+a=ށ�}xS�^3\����K�w3
��f8\, ����9��V�vp;_N��a;�`K��^��-��#P�r�fP��
��L;x���� ࡘ��Cǒ�g��*X}:�t��D?S����L[_����͜�n�F��1H����!�c�,�g;���?��<ߘ�%����z`�(\}z4�޳��Z#tڐ�Z�(��ԣ�]
 �}��`���'<�LG��L �&�'ϗ�7 )ͭ͜r���M܎�� OLZ��P��B�R ������.��9[��EqVp(���{��곞6m �Fq8[-�(1����n޽`�������0�W4�,�$���T�/d&a�����%ƒ�"�3��ө� �f�k�)��x6��⩽�	;1�ڟAϨ&�(�_�Z-I��HPbt��u��&�G���W��ӓ^�`�5)����{��l.�<�I�� ���lt����apB���:3P�A�ux5���e}/�����=��I ����'����+	-o��Ȱ��@Wi�y�*�K#eϧ�)�_53�zD78�[v!+�:����۠��AF�.d���*��G�?�/�x���-*$:�?� ޗ,�Q� i��I^>�����-)��j"�[�X��خ��6^D�۞?O6��2��*:WdO">��D��*x��KX�Ru����=��[�X�3� S�F���E�,h}�X�kxS.��9�q�M������*X�K���X��H�mc_P�x�����r��bjW�rKz�&�]���0&��4~	/!���@�uɏ��tf��"������d7�[�a�g N���@-�C�Tn�14�BV���L�AO�0���pQ����23�D������Y�ѡE�{x���w�:�.l���kU���DI&�Z*��we�h�9�w���
tV�1���Sؓ>P���.��@(��:ܴ[�o����fƩM:�ů�\
�F�tW5�[,�BΜ�P#=����l�#�2�VS���I�*`�J8�
8ɞs�+�<�Ocd�=9ӊ+QFL{uP���#˙Vs���c'�a8��:��iS%k���~��9����p�'s�#�ڼ��F.-V���!���5ilTL�j0l���a
MIv�.�����v���:#Z�K�o�9�B�E��B��V���ʴo��+`fN�Q��)�$n���?#?�������S��%�ۨk�:;�֎k�ˣ���*��5Ӑ.��b��%�Zr
��ȸt�P���c_�&��a�>!H���8
O8͉������~�iv ͪvƍsK,���:O���&����3g]���[)�5�=�_����n��Pш�Y#xEKv�y3��c`'��,�o\O����}9Bc<�N>X�ƕ
6�*�JƦ\,4u��>COp���m�&���o���m<P�Y72%y�{�?��0�j����^K��ٝ0:)�s�M��4F��Up����x�2I�,�q���
XO�HE�"�F�I%�RK뤁|F�»j�n�{����k'j?�=S�����kॴ�����wW�u����P�\���P�ڷ������F>��R3ͳ�D�~�[};ce���c�{���_� �{/����'PH�ɫ�yK�wCU��������oT>3 �:�kHT��yĸ3#� ���@��QJt�>z2����4k�e��=44�,m�'�CY��4.���e��қ:(ˠ��,ϣ�P��z7�}�6DG��bY�ƍ��е�dC�#)>��e`![�5��R�.v��2_��!�I��>�6R�Q�N�;#+��\�9e.�z�2���o1AĬ�P-���f��b�^ᨗZzܞ{�d��>����u_	�D�L��\Xz5�icJU�ߦ�E�[�j�B�^�����>�����"��-�o$/"b�p��^Gϋ�f��m�$*�X�_d<�Hp��l.HYg�W�@�}�Z�X�<�EO�,� u��/k[��nk�,�ϊ�e�l���
���c���cZ���v����G�{4w��(.��B�9��}�ܟ��ȴڗ�t�:��ʆ��;TM�v�J'�)��Zϻͩ��UTQ�F�������G2�X��g�'�����Y�n[�
����'�4$2hX���~�ѥ� U�ͰB�g��z�yN���
~ԋ>BE�SF���*����%��,N��k7���#N0ú��M�d �;F<4��G�_4���m�Kh�:�����~�D�.k��{H�����%�qq+�u�%
q����>�x���������ּ8��KK�Η".d,*#A#�w	��x�.���P���(8�^��/7���2�!�=h���W/�NД���/�2�`U������h����΀���]��(��/ud�<+tpՑWwG=k�}Pm9�z	��t��751D��:��)����}�A{���a�4�����Z�E�6�;"�֍\O���@6�C�L�F1���� U�5ܣSj�a���W���_3�MZ�V�1<���P�@9Q��G��D�L�w��Q�������5m���U���^"��;s:{N�aI�ڝ�e��|\ޕ�´$�y�^ׂ�d����Rf��Y��6Xĉ��c��y��3PU2��j-s���]���#���#�s�ԩ_M��#�^Z�=}�����s	$��s�Zr�426>��ۨkrJ�GUMv�͕��L�C:KG��=���+:���rT�t�|0j��q�$�+�qK�'H���"�Œ��l���G)�Lv�"��qe[�l�Q�@�A*�X�H �[�cU��Se�Ō���7X'v�d3�!�Gs�OA��`S�u��/�
,��)9*_�{���]x��G���Z��Q�������v,)��7W���i|��q��J��E2�u�,!%�,�)�h��f`ǃ����L� ֲR�Z�z��qT`�����B�~�o���"�*(/h)7E�Ly�~�[���T$8��J�6D�>���� �W8U����q�N����K[��)�{F�=�z9>�1��Y3��+6�7�x�ԍC���i(w�FW����~�#E�f$�atH�~�4�R�^�L<�q��{����Z͸�ħ^�@ς�=pGMq��|��)�ͪ�`��'��J��U�m�E�[?~=�ؘ��;��y{��p#֊Sʟ�Հ�A$�R�F�+�N��:��~�mQ3��i�
��(F̓��ܩPwLJ�Wzo^�3�Ď/9���ЬcEY@����8F߶�$zӓ�i����I�w��	h���s)~�%��#Z�F�ѧ�[/4�MDi�ޯ
�T��@s����`q���(��mi�JvXш�7�#A)��ς'�3�Y9�S��|a���E�J�	��Yd���/mv��t^Y0���>+IL$f�;�^��]R���\���h���F���d���c��L�3�j8{��n0ސKp6IZA�
��i���/� }�ƀ�y�� P��Ϊ�����q��Ka3����U��y|��R��L�Z�K��n�R�|cu�V�ǰ�ن=[s`w9
�jSQ]�ܶ�>tH�p_�c^�>�/gEϟ��"�k���p��nw���:�@�G5	R;3��0\U`η��1�;I���$��IL}�e;	��ļT&pBV,��� jVF�xV>6<cT��P�/�ݖC���b�����cAKQg�M���o{�/;�ʴ'Uˍ����Z��Z/��qf,�;m�ˤ��}�z����y	��L#��fr'P���XH��el�hk�b�c�q���!e�D�h���$��AV�ʔz�{
/�U�AE#%h�E6V���+*����=]w Rtlg��!�UJ����$s�d���[S�i�Q,Jv�\�9ɨ���;��1�5�ܭd(y�l�-�[���m�ӑ�[��ᐤ?6��ʉg�6�U������!�ǣ��R�7�}��X��!{��V��=Ғ�@
���㛖��2u�X$w3vڻ����uo:�d^��Z�z�?�ݲ���u���	���(Y��&�Oy q�\|q�����1�$����|�-������Ӟի��>��J�b?��>����Ot��^࿝�0
�<��5ƉJyK�~޾X���	�,���L����<��2��;��u�ղ4�u	A/sl�>���"6)�Oݻ������禘][r��֜!ȇq�Tpq4�5ܴ�/B�^#���,[<lT:#��b�VU�G8J?+�'k|�Z���4�2�����J����qw� �9��~@���=���o}m���P��}�rp���;v>���S_a�i���^�BAև�,��G7�;�����&���}&
*+>��\ܣ����Ϻ�c�%:�2��@9���x�Ã�� LS�Wrl���PP����.��A ��e��Vm^�?wѤ ��vCS���/����4K��ڣ�B�z���I%�D����&��ZR�Lr�+�:B�7|��D�6�`�?l�-!�'�ۚSH��ι9�OT�0Ɋ�]�����6��i�U�U��\&�
p*�p����$����=�2�C�&8��X<��@�I����Q�Neh�<�X�5;�(���B�Z���3e���܂R}ή�p��ֿ�y��(g�!�K�\,��
�E��c��l\�xU�6ocP����Wj~��@�$�Ȁ7�Lp0 &�b�sו�'�BDE���	�Bܦl-~��"���:�]��L d��0_8��������&�p�x8�ў|]�p�t�f:�Ef����&@� yf��F,���|S��:�Ls�q���X����Qdu�1����� ���gj7	�e�I�R�rW�<Ipd�*���y��˴G��S^D֘��wn��:Q�|�3���B�_Ӟ�o���"��l_�=2�0Nܫ�%)�b�z�K��R�g�Z��U���!��j��	l�> ���y���P�5h:~�&���ybc��n3��D�̓���h�d����\O�<��!��ݤ��r$_���B�0_ȧ��ߡ?�0��Gk��n�R=����m]vn,\��*,�)�/ȇ,;�z�<M�ni�=��M�Ϗu� ����lC'���2���|γ�L�F��I�Be�!S�f� 3�&��a���<ʥC�y�H��>K���xF!v�
5}��<�����	���J�ٷ/�F�˾ɑ�����Q�^��6����9݆� ����x~/}~�zJ�/H����`�/V��J�n�q_������fb�߹}��mg1��M;J������r�(#/�	1:1ݸ<���;](5�1b&���8���nC�>wЂ�J��rxK�'�EВ�������1ƗN^s�(~�{L���}�>s	}J����!��[l���܇�Uag�T�TI1U��(	�# ��&���'���Y0��5<e����k�����r�Y�:(~�«��t�n�����#�2�{���ؤ�;nqPn�8_��������:xxJ��d�#�G����4��V�| /05�o���wk�c��o��\)�$d�U�E��:m�hG���ύM"a3��ls�*�(|���^7gP�}-���d�ǿt��{�/���"�_ؑ:yt�f#Z\)�r�`�	6�j~�	w���[�oIo#��D�����7�u�5�soCJރ�2o(冦�KQ?9�js�닠Q���5�������a�ߘ�vn���Sڕ���q���G��Y��<j0��L5��q'�ܐI�k|-j)�^X�@���#q!!i��KU;99�b;: 伨o�Ӏ�mZ0�7������l�T��Y���z>,�~�������G@ts�=Dۏ<Jz���#���_o�Vs�I5�A�ᶺr��qX����6b$h�9�&��ck�_=4r�#2"��~��ޠA�z^#���m���a�h�eŪ�D���
�v�qe����sF�?�Y��k��	�\7����-9 H8�9��#ê3����vWs�6TI�LKk�
<-A/F���	�5)�<��@9�sp��� bՐ8�X^�
�Z�p�ӵ��r1�W�)��&�$>����UX[![�z��d|YQ�K���w����X�f�����|�m{����4��2^z���w�>�
��A�+��m��3K�k�I���g���볓.�j���~���߲O��U��+&�Z�h�-�P{CO����RgR��z(�@�Oa���E����Y�i/D#���'5Q�3<�K�_w/���n�6/v�E=ڶ6�ʩ�y��$C ��Ai9����͢�2K����(^��nX@�'t+\DQ�熧(�{�zp+,��Kh�"b�  �q�� �1���x\K�Dk����m�p���%X�b�5�7�+�� �2r��܅�Ç�J ̗�6�is��U2}8&����]�{d��-p��FCK��j�<�LږR��󣱽8��~�i��źS��S�F���]t��nP	CN�+�CJ���+��X�M�4��tY}�i�]�=���°�K��*�ث���(���\<7,�sމk�q|�5N	1Ϙ��b�O��C_�ꐻ�A4Ph�f1�����י@�ԕ$��H"�� �x�����SLa?��h}� ���WC���Ӷ����A+b�SE#�e�kyw|��W�T�S=�o~X+R�	���pe����v��v-c?�>�MPHx0T��8�r1�O?�~��h��@��z('��v֠H��Z�vS޺�v���u�X_��.չJKI)��9%Nz`B��;�V�A�� ��Ƙ�/��C�/�UKO�w�����P��0�{�y���Պ�O|X�.H�����/o�-,
M�o�T� �3<��L��v竈٩x����7���!-l�yB�)��w��ϱ3�������ݴ���,���\���P�:�����!F��!�����ۊ'����w��Z:��N�{,� �'.�q$1T��xk�\e�����Z:ũ3>I��|��d��G�]�/�N2B��B$�rr����(�w��=8cx��&�`�	�Tez��X��C��Љƌ}o�tc^�W�K���(D���J�K��V�2�L�I%K��HP�խ��cܬ�e2p���h7�x\=��.��� �����NH��>ϊ����_ ?tY|hF t������̗��(0Bބ�6[¥ƱE�8�~���4v�����z��9�)�.����!>q�P��^���% ɻ%%�%�"$�n'>+!�<��lB��d�f-�N�P���l��I>��([��Å�V��OK��.t/6w�XD}{5�i�����$�cZ���u��H`J�T��O�
R/L�o��;����՜�g�w@h�&�FJP㨶�"�38
�e�4eT6�����d7��E�z��V6�7���5�Fݱ!Gd�c����[�1��0l��p���G��:F!��jU,�&�#+W?P�$����q�$ꉫ���������b|��~��&�,JDäƺ�O��D�VC��3~k�A��F�>�&Y4�#y�}A�9}�<9b2�r�Z��N��zG�*T���RܸM���G��,i���	!�V�US�9������#��i>V�3���6	IsFhY�1DP%��i�ZBc+( θa*�\��j�;�Poc��\X�w_R�yi툹��A� ��i�bT��,�#C3!|3 -A����b0o
��j�`�D�y%<�([�w`vJ�!w>�(��Q���s�"�s]x����?���Rk%.3 \z8>���JIھ�}��dsd�2uo_�����ѕ�*WV2Я����^��s����S���:��y��8�����H6������̙@�(#L���g?
���r�I���)T���lb��}1��l�.��V{�!��s�tA��sV/<�Ad�'���V�H_ڈ�"3��L6��g:]3%lO`&���*�<�J�^��wW�߶�P�W�er����+��h���o
���������x6!R>
�Wo8蝢6('u��F�W���P�`��@���Q���MA��R�|����isS��-[Y��v�5g�?�z9�g.�@+{��~�dI ���Y�c-��B-�Q'��5�f�T���8]s�o���{�%��3�C�Dq<B1z,����:d�;&��&$\����0k |���E�L��]���7WH����H���4�=����L��EK�0ݣ��lm�=�bv�\��)b�@������,�F��$��y���*W�O����5Yf&s/�����4>�Ȼ(%���C����;ٳ.�Z�XB�B��w�(N���cA�'��v��'�vl�AQ�RrKOk#H�ᏇV��w�VO*|w�9HLݡ�@���.��a`L�
[T�����!�KbQ/IO�A�kOv�8�Ӊ�렐?�<G���Y�)��pW>R�L�7�,uZ>v�$���\l�ՏV�Y�ՠT5�}��zy�$�]��&XE�H=��!�l�X��7�o�})�e}�PhTB�.i�2�,5nr�J���;7~wS����{���Gnf�^V���cu�z@�~�Ϻ\6sd�s$!�-���0�HX������V�R�Ю�F�G%� ��kZ��nY
��5��/ļ����1��,�+Ζ'+�
]�x���%~;�9�r�bR5-]��~h�� ����$V�(�f�^�{q�����/�}�$���^n�<�xD;�oqT\�>��3ݵ�S<<$�u�FƯi'w�i��^�����W�_���Q�}��u�N�r�I4}�A�-���l�Y;e鎍���r�Ɛ�T�C��Ad!MP�����rCAu��Ô�L6K�<���5�l��^O�z�m��.0h)D@�HTl0+:tϖ"G��!]�h.�����6	�~ᑬm�}}�]jp���FP)��uMb���FfzE���V�#S)v$Ӌ�V����kr�Ѳk����>E�ѭ[��]͋�Tp?�Tn�4����C�eHj�ճ�4x�>!�����nj/_W`vf3{��d3;?����|�j�3w�s��!ⱞ�DT1�U�._ǃ�4x��^%;�A���~U�n
�0�p��揱�R8�~Ѡ�W�%:X>�P����:O ���,�[\Se�͡u!r�����n�g�麕�i������+O����Epg�e��/��E��`�����?����t��K:�8��I~*��Ų\�Rt�I{yeF	θ������e��.;���V{�3E9-x�{���Ɍx�'5�#q��o�椴'��^r����tI~�*����t`�U��UN��/,۹U�<�ض��c��8q�kW/).�C7��|a*�:�0��� �YQC8g˽-!nL��,�W:�։��G�ޭמ��)�@ �E� �ťܔ�P���7��a]B�V�Ťz��˳Z� n��:�4��������)C� ��iP�"uұ��]S�>!�����{s\�xb5��g���Q�C=��</a�r~f�0q)���L+m�1)��{7`D �f-蹲.g.�|Վ
�N��&��5�,���"���3@ߝ��[��y�r���9����+@2�xd�(�qcd���=Gp�^=�1�t����;�j,D$�c�s��H�I�!��Ĵ��s��q�� 3���;*�,ֺ	���^.N�&tfg\7|��/�kM,d.�4 ��}^F=��8b����o>�o�o�54v�%8��\��%
��U�G�X8`]�I0ȹ���q�+ƪ���-��:�22ɢ|�+��C�N㵬�@F�J�� =r�K雘i��)�΀3�[t"��4�'����f����>�s�)�(�i������yB�[Z��ٕƔ���;�d�Y)���6qD��^2��,�cFE��o@�3�<fԺ{x��>�kR���{��{��L����="Rg?���6��i�7�^~��i�I�a^Q.~=�$i�����\V�\p�g���*(}Z��\bt�mT0�n۠���
�"sO����^I��J��� Jf��6S��ݲ��� ���9#/G'/�{sR�������j�I�����5;F�_h"�畅w\d�@&�#\' x��|��1�i��V� )ۓ��h��&(��Eq(�D�u�ل��س������j���Bh�]�`2ޛ @ ��a�l(�� I �[i�[5>|zk�a0DL8���/�/v���/��3��|{e���-MTp���2������"��־�˘4J�������Acj_;�4��;>���"���M8�S�P������Ҟ�c_#,d��4&�!��񌠯��7	���2�j�w����W!������նwHxr��J7w���[��-VE�u��s�=$i+>A�d�Gpgs=�,�L��JQ�2	R���}+����T��������!��"�Y��/�(-!y�r�5L���%r�&��BCr�����'>�yX�b�'`���Ÿ![�������� K���ulS��߸�ݫ7��pt"*�zN����ɞ\�S~�v�����l�J!d�Q�֔�;i��½M����hK�ۺ=���p}Ӕ��0�a�@�YC���#�cy����ͤ���)�_|�3 wTg�?Np�=OP�T0��,B����g�^����	�_�\o���S7���1cC
��cm�Kʇ��'�O�h���C���y��xz���{�7z�m�6v\h��yM4�y����[K��9�c](	���'ѵ�Ch�&��*N�ؒ�b�H5�B�Oie���%�|K�����?ۆl��E�*���|��ؓ��'�L�P[���l�>�!���*��>&��������Y���A�W>������e�_���|žm|��=�E��ުs�c��^�$]sp��g,�ܾՉm�(8b�r˂s��x���@���к`3j�1�\UΨ[��Š�vܲ��B�y�鑜�4�����q+�R�nK^F@X�-�W�*�%��%�{������	/�ε97b��Zz�)掭i5��D�|�~(gX>.Y�|��l�ӓ���7�N�Ca�r�8�U<��"��&��F��~µ"q���zP���B�]�~:׾�(�"�!&�c#���=p��~sK]�������:o�j�r�G���bm��T'��MǴ"	x�Ű�	?49�E��1?ak�%~�0f�^��Q��R��"
8��)˱�������s����5��}��xt��?�Y�A�D��y������El�&��ە�l IL[�q�k�X�]�K��^�Wַ*$(q�3�(j,��F�J��KGظk�r]�x��ǭ��d%�|�,���|!����;���qi���HimOY�Gq�i�,�w� !�A���������411R� a
��`�l�a;�r�bX�k�)��VеO���{�N]���y�������-t���S!<� P�c��pT=�_\�Y�i�OH�~&�2@Ӹo������d$i���ѵo2��M���*�t��A��	�}yMK6
T�]
���i��/�nZ�(��-b)�����.쀠�C��j Q�O�f�<�"R�Fa;(D0.hH��F۾��d�\�k�N�覥4��x�����~�y��dC$��J�3]R���7ʥ�j��|�
<L�U3\MG���
���BF�A̡ܷ������'Ė�ƪ���Pz�)Ā�>�;$@�frd�.O��Jʕ#4�( ���|�\c�5P/2f�Üڎ�z$D�*�̋�9پ	1� �vҪ�B��EE��p��o'�5�2,'݈��E(��p|r�)JV�ɯ���sD��Y@ہ�����G��}ozo9�ڊ�Ьp�%֟����}|��*��?�sj'�ms !O>MI�(�ѵ�:���@[����V�bN�@��#
~���U�7��[st5�p������<���Iݲ���ݝ暬ڰ���=��۩IZ����#c�L��\N9z�K��FQ<�	�Q�����y�&]���d�����1��\/���^���^E�,l$��k?ݬB1���eg*�i�S���ѓ���-M,�]�	�%����]�M5�w�>N	xJ����剜p��-�=�K�"
��������?H���䁗��y��}Z:O��AM�Yv�����"�O2N��<�@���즺t񐚂V�I�Z�q���Rn���5�.�>���%��44�
�=��_��Ǩs�gU�ğ��ׯ�}�C�4�	�l��7&WZhCm��/�v4��<(<�$-��Bmq_��P���Wi���y?�����^�Y}qPhz;	dj,�T��Re`�"7���˚U"�x�����J\h�z���N�=��A7'vt���7yMp��e� =>�����g#t<�B3c��2�\�&�%�@��{���
���� ��o=,#9�>�&$�癙����Do�E�,�$f@%�)5J�ߍ{K p�N�N+$#�5?[�*=ҵ�7�gSW����˟��	|t|�%�˯B,��Wu�:�m��#�� �n�#��`�����O�1E�Kz=�-���ǝ��B7O��<������z�Ӡ�VmPT��b9�����rH�j�,�}i{���Ȃ���f�q<TO���[�#u ���0i'�_B�h���c�:��壯N��aƹ&����1��L��\ZB8��� beCN��ue�ۏee�Ԕ$o�n�ؠ(�X��@��m0Z�v��i �7�g���a��?�,I����������U�~���]A�伮u�B��y�[&�£�G�K�ސ�����!�$�����v�,E
�/x���(�v����g�ψ����H	X�l}�aiz�k���4,�[�vJ�.�ƹ�p��(�� ؎Գ�%�=����}K��F�}�5!b��� #����6qF�� Y�Y|��*`F�X�wF+W|`p�\�0˰Vڞ/��F�ֶJ�f�M�GNR*� ����
؃�鶖��U�m��]{%��O�A侉{�f#����в��9��b�&�b�Nq����7c��P��(�:F���*>v�\�]o�o����!�����ә�K�ޡ.�wp���G~�%i�Os�g2�U�ƫ׾�#�Lu�w��~�8�V`=k����H�B뼤J��R��������bR>���`��ۉ�5S�د������7����(��Pװ�،ge8��7nbw���-�;�(��� y�Q�nӞw4k_B�y�*��B�ϩ��J�!�9C�@#�s]�5e�0q���Jt��\tB|(y��7�d���� ��R�t�)z�T��g�����){�Kuݹ�"��g��!���i����Ɗ�u�����Ԕ�dǦ�����y�Z��Nw���y�,|�ӊ�E9b��ɲ䘆 ��R����d�Ն*^���k:�@�^��T&h�}9ZD��aݍ�΀BIk�
huY	IP���UC������s��Ww��Vؓc��Q5�l|L��$3к�B��?��ǥ8;�J����E�@��U1�f�?� }W�p�n �M�i���]�Sl)�3���k�/$�����{�F�KC�Y�H=�=���0~o����n��z��G@f1m]�nK}-kb;ۖ�j.��K���oݳ�z�����A}dP^��xܡ%�я�0��Zt.C)����}Ƞ��3<٭��x��!�/n��
COG�����թ��r
#���h�(�+1�)[��sQ�H �CS���2��`�{oA�]���y�����:���M�{��*��BI��<��Gv��{��ѠQ^��@86�Q�)��揶�I��h��o�+�P0ְZ���:t�|�/���ZVk�nY���kq��Ro�響���W��WhЉz���C'�72�k�zJ���L("��;�K�����Աz�̤����q}DO�I H��Һㄏmru)�MN���NQS$l&�3�o��ĩD ���uN�)pӑ�u��@��S���>�r�x#���-P
"�Kʪ�߯���Ţ�q���5�@��:�@��z�mm�g��Ս}+�����M�C:�~��k�ڭ��$��ewko���%�rB�xD�P�`s��YM����C���R:�jE4��ǟ�+�ZC���RZ{����4aƇ#}��.G���6��+�tW����h�ک����L3]�sq%��iۜ��1_�e'k�Z��m7i3d�*�g�9�\h�j ,���G��-����g-��R�T16kI��8�w}�7�^�({Mc�R�p�J�`�j�#�(˖]�9�L���$�bK��8a�J�P���i��#)?H��U���^�U�v��s}��tz��/t� [f�T��H�Q�qՉ�&���1��X���B��9U�N�~)F�9�Y�b�y�t�?��ZG�����9�is���τ�|�t�?�/�๽�̓1l��0Յ���[uq��f���������H���6��j��ص����,����۳���I)n��B��P�������n�Ւ ��Q9��4cx�4��W�W���!����!�ҿ�iL=;���F�W�)�|����N|a-����w8���] �9\c=�J"f�ŕ֡i73��B����Lu��6)�y���P�����AD�AU�u��ts�U�aŀ�?ޖ�Ynw_C$1;z�`��������|��`�n���� �l\b�o� �����yb�n��0^����������e��h�����{��/b��q�o?�V�e�����B�C+��?������M3g)yo�m�lok5��lTvc���끆�N�.�=Ytbγ_/� ��s����ъ_y�}�b�H�M�ϥf�C�f*w����oZn|`3����I����tcx���u��#�^��������B�^e(�X�4��J..�i���ֺ)�d7L�:�'/8��e��8@TZ�t���V���E�=iz�y��1����W��2����:�H=���|O)��[��I��L������m��;X�Ϋ�"�|n�,�wJ�dX>�gV�\~^�=�a޽>TЀ���`x���{/
��ZB��\�����ՖNQ]xs 2�q����!HD�g8i�7ϣ�������Qjn���c0MXV��g��G��

�T��6���C;�i�ĩ���ڲh�\$i!*�.j�{H�jV��Q���b�J�):��3*�f��OO2��!ȇɂ����H�xLdءؒ*C�3m\��S�f����q�}̜�`F�����:�ց2��6agL�M�ڜ9���
���4K�
2z!;��z�)�i^d�쟾�İT����6͆���7�$��{'�����l}N����t���z���g̒(�Ҟu�k�[}�I�!��z�z.,$�Y@�%.�?��S*E[�!�gZS�i�Aʨ����+��";���	����4���N���?�tJI�������s�va������	-K��J��k�?���5�5����K00}J�Ή���[K�G��br��Cr*ɇfx�n,�1G�'��5=�ƾ��,��"q��N�ptHZ���2��
���v�o`E���{��o_�$n�6*)AF�!|�^H�^QX�ن����K|SK�`���2��T�P������ͯ�O�%'z�2{�*kf�[p�*nF�L��m;�XG�N�6�@S�X��]�0���ش��JK��ܞ��a��Vk<]����[$��e�HA��^hsbD�Э�ݒe͜n�����q!l���V&��<��~2f0_m��T_i?�|�G�.�X+T�>$R�Y����Ygj���מ���2�x��,�-�Z�&jGC�
��Y\��}�g��1m�ܠⶴ���O����9��p��@���pڥג�a!�2��\«���<u���l������Z���m�r!W"�ꀸ�-.��3K�d&�ʳ|uK64i���Q�F[���z��Y��{W�3��
=/â��ǃ(����nJ�D�c8gKf�Tb�L˼��J�z��;fc��؆1��P����*c�KЊ�8��fJ˂|�OV����M*:�!	� _K�pm�Շ��(|��b�EF2aUT�[��zf׵���a*�6��͝�L#����3݅<w�
!����v�Jу4A/������ʆ�=���T��1���E�U��w�.6��5?�-�z]�GJ?"n�5D|� �����MZե�T��` ���l�%gOI�h]У��m�bl�� �?�3ͨ�7$�0e��$鿰z%�C��H+��\s_\Z�3�A5S������4	դ�h��r�a��2�N�s@PPL���5��������Ў�i	*;���ո��GR� �)�\��-�c]�˻�,�ۆl��T7��w|;i�����if�����<_�5x�m��Y�Ip$/tɑ�z�-���_b�r1i�;�DZ��&c�=(��?-� ?J����V*tkJދ���y[�^���w�Ok��7Q���z{4�u�KN��-M����ӎgL\1qyF����J:�O2ZH�;(j'�o������r��,%�!1��f�i���;�'M�b6|H?����l��SC�����>���'V�+�cy^?Lɘ�#��)1�Ez��&=�8��5MG�G�`zN�#!��� � �q�f�֐-����Q��=Q5�_ޔ5Ӱi��v�Aw�u�Թ��D4�1�������Ȱ�9���w �1���l	�:	�ᬶb��#[�����y�%�%�����+��\�,7�F�y0�����Z��i��Nɮ���=@���5BH��~T(܂\�%���,��5��)�F!�^�O3�����	�"��z*��1t����%��"�b�t�k[
���y�Pz���>w*��Q��B�  �q�Jb�cnX�RS ����b�=A�1�L|e��T�ಠ!��7��b;�A�"��0�a�@`Ɇ�$�HR]"�/	O���f�����G��#F�b7t3|�N{�OI�}W^)��y��^B�s10�1�������{+�eLR�
������IGm;�YZ��4}O K�Ҹ��1L����
}��Ģ�pqf���첚˂�-r(2�q�d�W�=Uv�o�T�um�J�4tuF��$��6k_k8��>_�9���{�
�T�Ȩ�������!@0z}����!���r��k�n�m?t�^�,�M>���Rg'-�5�y<t}�#��'m�,�R1w��'�T!6����Α�l��|Sp"�M��aɿ[�/����j���
�1?$�b��=�(�I��q?��%eM��K��.�-v�r]Tepr
p� k-��]j�X�x�c��I��4��bY�ؑ(����1�'�8mU(O�����O�#ң�\����1��)���V����V%.�DPG�zڡA�3�ȉ�,^���⩭�m ��3p"�U���ec�7Z�&Yt��s���������.���"�1!t,qs��][3BU��L_�j�ȩ��S�����&�(�/� H$N놺������Ư�=w�<���|����L�,�Ƅ����dğ-�-��"<�U�Uj�S��jן��0/x޷+a�G�%=���$��{z��]W/=p!{�yR��0����(�cq`ΌH��z%\1�+S���!~ɴ4�`������.F:�����@��������JR��{��34�'C+h��.�� �0A��U�K�YY�v%�-�@��mn��}K*�5;�O����ڞJ��JI�40Jk�Z�:�xpY��� E������*�'��,��G�'�zb�2C�����Q��� m��Y�"6�8���n�KU�C��op�Ӹ�`�[��A?�k��^�H�rw���m���9���Ad��Ԩ�!S��D���u���q�Iv�s�S�����
x��-&��,8v�%_(l�cծ�l9���C�1︟������߳e�9$�	t .ߗ�S�h7O���y��X�����'���͞t�x��/��i���q�)�y�+yщ͊k�K�I��?��K�ΊXX�McZ��gئ�$<����0�����r�Y�n�S �T�.L��8����I�"���w�ܩd�9N"��Q���J��B��P�b����Wt�� ��B��8��ɺV�Ƿ8Ԛ~Bud����|ie�N���k�?�R��d$ �������b�H��Y�#T$5,�,�PE&������a���V�1�y���e�	�5�� ��x�)8]�2��Kw�"���}�Ԉ����5�t��R��z���=�k��D�l94:t��i��XC�pv����^��N��k�ٙque��_nG:/���	|R�h�W&�i�+Ǐ�_0�uu슕ф� ���G͏G��RQ�Ђ[�nd�N�铃����ehi��������Re]�D�h$ܚȽ�ꋬ����Gd4!˧�XI��na@��fjo�̷��oq�HҒFָ�9κ��69�ij��4�B\�x���8٧��@����;H�����D:w{�ȧ_��DO n����<��� ���i�j��Rr{-i���r�p4��V���B�r[`x�ϥ
�hٶx�3mڧ�>Ձ��*8��T[�K+ D�J`�%��[�J�����_.�DH/�)l�o���f�����#Q���v�y�,78	y���U�Z����]��
z��1�ʡ�pD�h2`Z�BK��[Yۯ��5�%g�lf�7fY�t����&��=I����?WK0�(�_,K���Wmvg��h9i�\v��\~]e�ƅ����x1������56T����p�q�^[�;Wl�{��vٔz/��j��4�+*�Y뭊�.����WS��|`�Z-d����)"��ڗ������d�ݪq�x�^L0�.�Y\<r`VXR��ۊ@Cl����!�=H��aW1~/�
<ۊ춎�Hq�/"�v_��%.w�4'��o~�C*'?o��a���\v����q,�4�J�C��i߿�y�?�1�0��&����8��A+�UE���'�'�m�!#(���!��s�S��t_�'�>Ó��6���p>CI�Bu���$��s��ױ��!�`��O����E��- �J�Wx��>1�B�'h�#�)8��6�kȏq����{����@I�Ŕy�[AOZ��O�Cer>u7�R"
�4�K�Ml5�_�E�B�y�-M�n�yIN�6c���, ���yZ2�FR,��Ϲ�#JuB�ŕﭏ�</����g�c�L �I:�\D����)�h
k��íz�,����>Z�,�sb]8վ۳�����7x��MTw�dθ�����x��0؂��*���N�V�A���-P2X���]et�!U�E���҅,�[+ǐ�&�����e���:��%&��D�)��V*�&56F�!<���$����j���{����<�Ym����� �(���
�$��"o#��]� ]�Fp�ص�x��Dl�� %u�^��3bM�x�z�F��~7Ȋ�3�X"�.y��6��?f�R�l����󶶃�>r)�z��z��y�p0.s��=���ޗ�|#8�"y��Z<~����P��~{C*\�/�8��C%0�.���F����w�).�\�����?�|A/�9�!)P*a��q�8��ax����t�B[>QtIm�[�~�*U^\{��p��Ѹ䬪.SK]����R�	���RJ�*�48Q��`_!��8���^$@��j}�gc����Us��� ڷ>��������N�B7�Z�g���o�Ji֙�,�h�,�[\AFIg7wS3wV��aQ#��G�#ƙZ�`Y�Ξ
�I�C��"��\~����k�N��h}�-UB�9�:	�+�e� #$f�6�A�ٱ�t�S�I\��^���oD��B�[�8��߳6C�����@���>dJ�/j��R9��]�z�yg�}$O�D �ţ����\�q�������|���g�О�����m� U|��=��X��S���T��Ah%�����Y��3���D0.�<��KUg�@*3�LS���;F�\ ���-�|�$Ej�^$<�i,�3������(��kF\�?%�7/7BҎpO"�Og���;����|'�~�w��N�<$�!��l�OA�r&=h���n<���rGčb:������ӌA��A~�i��H-�
���ΐH,R78����I�<�q�>�!"���Gc���ճ�=ur�k?�F	�	=xL����	^�ʴG�0�z�{[����Aն?�4��'��ti�_uC�Q����K����y�ďs�f��aI�4�ޑ0��������en8s�5��/P%�\��V�ӝ���+t#_33+"�k�[��p=�V_�3inU�4R�~f�Q#ia&���7����w@7����8�[ ,j�
�Y������)��*��ˋ��9�]s�C��� wyVj�(=�����c"�nV�h��j#EJ�'�����W)�wQ�(g�_k�� A]�I�"�����>�j0�ֹc�A:Ӝ���kq�ݼ���;я������#t��=�Z����v�}��km��ƛ���ی���c��/KKIf#0>�ھg=�e���#&=��c�5��X�vHd�2eb��t[4�����&ų0zn����V�5���#�������ۧ\�͋�j�SK|��u3~�^�=F�F,�fIs
�<�
R���қu�\^��\�m�yL.{�şf��:]��X���_��hn�gp�ڀ�VL���s��7P�DN$��^��qd�������z^��ᎰgY)��� ��&��'lq�a"�Nt6�7d/�hj�7<Jl�2��t���ۖ�/T.����0���z�}i���]��Á���q�E���cdu�a�U-�H���3�x�]�Gg}�^2��R9���P����=h���co�w�W�:>aLHK(��D,�<Q�Z�����@<u \������G�̣S�O�[�8�����T���s���;U ����.dS��G�+a��\ �?�[-3���k�[Eoq�,(`��ͷ�����$��5�(�� ���V��m&[���}���,u/b��h��59N�`�����b?�m��Bq����G�CF4������u��a��G�c2��{�c�BF����<K��[䅛D_���팲��P�b%�R6E�E@�ʇ$Q�ū�&O�}Ĵħ$e�4�6�����=�^��f7�i:�$�_�NZ�v�%��l���;:����}ڝ���>�P8�T;��jN�a:�IA���l�>!��y1^���p�� ��OE=����\jk��.�sW��"�$����=�_��"j�q6y�y���k�I��b |��ql���%OAጂ��$�[��#b|��"�+��	��ܓ��p	|f�,�E�ӳq��
���Ejd$�cVJ�X߂ivJE$~ߪ3Qϔ�dJ�1� |�L3_�#2�a��jx��j��h�Y<�g�h����(�Q$ 2 ������=8R�ҕ�t�jr�n��K_5��a!��h�ݣͱ�?�'#=�C�Cw�׫�N+(�/G{���#�H
�UL�/��ŵ�Dπ Gq?���9��W��KL4t")�]���ab�l}�.D&n��b'E�-Oր��*�)}z+�9��챙���f�9+�CT���hp�<@��R��n�t���Z}����.�Pp�LtQ{��{���`:��x��{��}��i�M<�&w�7�&��s� N@I��p&����/��E�/(�Bt�P��r�"Фd�`XOU(M�4ptrS��D���=̭wTj$Mdz
�X�� j��B����~�������D[x,�p+\<��'�M��>���O��q��i�w�掝�7��C��$P%�ߵ�r��*�kذ1�0�1�۸�^V� �t�5߶��鼊��UL讑ЉζW�Jz<шLn1]��ru/@F�X��S�~�x�	4�����8�*ϲ��@��4d,�h�'b�V&��Y|��(Ft�%�x��Sl��ϐw���<[c�Ͻ�瘝�����/m��r������7&��vD��+��A�Q*����R�T=
Y�T�~�h�F��0��CѢp�Ӑ�Z��Yn���� �]�.�d6�P,��E|�5�T�ڠ�0r���1��Q2Q ���Ê�Y�@�����==cĔ�u�qH� ���Q9�����y��;�_�i=�q�ZB�����\���S)�b=���z�Υ�'��$�����OXh�����r�ґ�Z�S�p��fx3Z��P�!����H��H2��d&)8p@/`#z��?�� �&{ӦN'ìa��d�D�)}��qݏ�O���nx�9���Sɣ��D��a���_��N�DU������� G4
�~��6\,�J��y�sH44�[�]�$%ÉI�͏ȡ�sU�PѨ|.8�⑨����X�$�����Ȗ�%k%��ҋcDۗ����c�So�C�j�~�������+��wƃ 7��G��<+��3�%$(u�=9|����NC�y/����� �>�U˝?��o&d���0��ˆ��0��4­I"ǯ|��q�#����w��(��|�JP��������_���C�{H��M��	%3I%S��B���	:d�5�io�襸ff�	�>\�ޝ"Ҏ;"D^nv�?��_��\��1��: ��I���u;mqD.M�D9�LUY��Y��m��)Nr�a!��#@���,�JNS�C}TGeD�1��sQw�A��pB7�<�诙�&�o����V�r1+b6%�s ���N\� ���k׽`���l��P(��v��݊�^�X/>�OE uub`���˰{��6vS]ؒ���b��UO�
���+��P�Y:)�thT��(J�b�	�=�
B� y��M&rMc,Ь�#���??�>_3���⃑��4^s�J��ӹD=��H_Ve�MS���ӭ���S�wN)H	�`����~=�w�jFGO�ϳL0_�� ����g���Z��/'GJ�G���&)���g�;��ȩی�%��.s��h�N&�v
v�Q��A,�dS&/�� ��EG���tn�pI ?��Û�k3�:�޶Ӥ�@� �xDL�Y��}ť������"Q�u>�z{�3���K�@d��x`��}s��2�+��p�D��l��ԗ��_�4�򅧺$ K�7$��I'����B(%3��Os�3��j�w/ ��&&e�D9(��:�ྐྵ-����u����y��Le���c�Jw(�8X��y�m��<��	�9@.��eJTw�c,V�yae��&(�'���-q8�dp�x�$<��4�����',��W}h�2���TƁD�{��"m��w�C�.����T����ũ�V�3���-TZ��1=�a6O�Xk 	�V�/漛K��d��b���(k/�)da���?7�j�"a�Ưw���n�i�+rl�H��c�C��Y�E�Q��D�N5�r�)�`�C��=��%���]	�Q���N�s	q� ���b�\�6 �M�t_���&R�İfLq��n��L	���+چ'�Z�ς|�T���DU�S���	'�| M^�FLz�Xk�@�.3��F��ᆰ�Ǩ���jXIGS�юl_T�	��jV�!*��2�\!G�#Rlaᨂcx1,q�*g�bP��m;ܓ�3��ɉ ^�(��e[�ZT[��Z�D	�}���x����e�p�����r9�`j����RpyZ�LaSF�([D���Zs��P����Vט�!M�
�u�����E�`X8�P�)�B3���\`�?&��|l&��̓����3���� B$ɔ����k��[�?�c�����
���4El��E����:���������u(yR��-!�)gyA�#jd��ߵ��m#�[�91��F&�[5��x,�:K!h�NE̈:��a�W�8�7���2ɥ����6���~(b���D7H,�l�����Ĥ�x��)|��&ǡ�[��G�%`�	�!!{[o@j�m��W�]�.�E!7N�ܗ�')�d)݈��e�l���N�K�:;���εzF7h��9�XLn~�PAqj,��1��J�wAގ8�K^IB�W�iU:˒��RMm۽�QԈ$�O%H��l�e�ww�s+	0�w۔dS��d�U o"��U(�?I��^4���J������m2уp.Ω��"��U�z����v�\�&��jc���v6��7��P�6d6>:�JV��؄��� ��hЅUt�6�Z��f�ӸB�!�w�2����gZ>�M*�~�������y�n3P;���a�w��Gv�ۧ�TH��]���m�$�B؁)��P lo�VwP{q�)jM钕���4S�j;�Цd8ѣ+�[f��˗t�����f|CҤ3�������:.��j��7��E|��N	�8!��33p��#��n��;=['�W!j<q�&�!�:�����\�TeR��"u�����}3��wZU ����e�����A��\��aL��k�`�]X�@>Jhׇ���ID�m�\�а�h���|P���a����˓�60���T�����=��Y�.�2�6�`)���;}RdY�_��� H�(��3Af�>�橬�cJHU��ʁ��f�A$S�͡Ρ��!h}����h�v!��W_��x�gv��#����,?�k�]�/0T���!*_��?|�5dp�����H�c=�1(^�VFO:Q�i�i����+H����_&�����:�Z#d�@i$B�śܱt1T���Ա���[�J{�N�m��^�0_��("�d�g����	kSV(r�%-M��m���~����_�->��k��N���Mƭ�[w�U�� �#2<B;�u?=�yf�����e��ՙ�7�J�<2��B�u���r�*ڏ���V��`�] l�k�n~�u���f.�郸:Y�
j�bUkՁ�~v�m��>���e!���vp; ��1O%N�������v1N�g��B�QR����,��ER~{Ң��p1>禉���D��+��s�J�'P��~�R����������)����}���t�ӏ��gV��ٮ��3�0����ų���!S��n|�̽h�w��1=d�<��ti�]�T���Z��U'k��~�Ep8{1d{���*�-Y�􌨶\Y�{�}�?!�$CA3��!��9%���p#[�֮C��wCj�B맽O�4���A;y��h2-�Nf֒$G�`���eȥ;�h���v2%����IRS�����~g?�Sv�m&�	0fXģ�E�+�@�~��a�u�b�ƅ�"�b����piK�3�kUn��5�G�dJ��&�h���2��TA\z"�o��
��D*�Ȇ+�OJ/sx��?*:1�?��w�dĄ�j�)�.Izu�4�6G��io�n*���<�6$!��{���;=���$��(=�v���0H��1@Fv�dT���)n��`.��ÃG���f\��G H��a0 ����680��c�S�-����Ԍ�0^����\�jl��,eQi|�5/�*׍��0u�k��nD�Zi�n0�o�{?��+��˪�WU��7u��Dl3R����ѹ��~,��)����0mW��o98,F�(f˼+~��&9��ò0�8�`�U��M�i:u������>�?c:L�ov5k���=:(�x�����������_�pf�ؐ�+{P��6N�NǛh��^Pωs�uY�$��`tu�y��h���'���##c�*K����	{J`����*����H��.��'\��Vn��`��&ˈ�[�/�T�Y�|tU��b��\:���T��j��0��y!�������f o���nG�0����PV��g�v�4��N� ����^�Fw�c|y-��/���t0��rbKD�=����i_�]�t��]����B���w޿>X�¾G�p,C��1�ZK�*��.�D�O6�H��?�g��P�$��h*rI����P�q�ZҲ�x9ӌr�=W��y�!����_��7���(a�`�oS"{8����c���(��l�Oz[��Ԃ��߈�ǿ�WT���ڢ�~� �	dp��3=����|]ISч���S�G6��"��o �6w@�[l^}�����PG�6��V��4��ζKF�����!�a4&�f����2�J#o����c ]`�DN_2*�@���W=,��F���_�p��h�� *O@�3��U%�S��?�j��L=9�U�5u�L*�L��$'�k�I;;l�io�P�<?�s0�U�[:��}�,�(�1��n��@ͯ�p[��)
�dg����|�Xcy��R�N����	�����y'wg��,����)���M8� ��C�,��_���@�͵��pfHx��Vi��w��lA���F�8����.A�P�0Der�!?����EC�i�[$�~�f%�ģ�C�6,�.un���:�QA*�=��c��c!�>b�B�a1��4`'T
�Z��i�
�X_K3��o�?#����X?=��1uՏ�� �y�l8go���kqn����\\*F��4Ie��ӄʳ*e��ap��$�o��^��֏�
��:��ĩ~oj�Ϛ�F4�A�)�r��\)0��|� �bu�����=
څ�Q���O:�FA��}������A�z��X�9 ]����s-��G�g��+X�e;Dޜ��>���9�z�,G�����y�{� �Ut[��W�X�U���/�9�f�r���.l�ZN���;��s�7��������km�!=ˠ��Q���(Hb��@�u�\��4����S�vރ�"��?br��+��-p��� ��6�<���ڜ��hx{#<u�ʗs�����9X�js�4�Ht9j/��z,�������^�3������h�7�C��K�J�Z{���k�L���X�ne�W��r�"W�S5<�Á�||x)
��S9c(��(y�ќ 6�NF���K��z����o�)}S�+v�f�t���LѲw�*�*?��Ϛ�2r���b��C@N���۹[����:=�hj
M�wH�b&a��`����;TJ�+�i��~��2�nЊ ������R��WP�,�H��<��ַT{�w���e=�e�,NPII-D�_@������#vD�!6]Q�羆k��uSq�9׭��R�2,�i��
dB#��~c @\��w�k���Oy��]0��0�ڧ%R�KR�`W�D��V��Oӛ���p���L���o3@�G��$�x��4�
����*�_�9>J�d)^�!�Ɓ5D���e[��P�K��0>�!�ֱ�t4&�E��1��a[m������F	���-X��[����%��(��>��IB���%3jn(������F�
���HHm�1���;�3J�W��N$Џ\��!A�#
�[��Y�Y���{ю�Z������Q&BRr�l�r�k�G0�1�^1O_3G��O!��R[QFpr�*8ϐ����y�?��V��N8�^����K��LJ�_oó��ż�L�l��ˎ�=�I�C���-���Ύ�M`dm4M�Z��R�o��c/�Q��쒄��^���u��^R|j���Z ����R3�1s�BP#I������%��v���i�{_U�Z���<<vS�n�Ym�������`��D)�H�7P����"	^�{.�!�3j�Z ��ȩy�G�I(�T��G�T��h��a�:\=q)S�Uh�
YԊw�t�� A�����N8���m�XKH(�J\�M©��?��R��5A�N��Z��q`b"�S�U�&�_W �;{�v���[�b<:G%���}V��x9���:�7���c(���w���8o���H�\����h���WXB-*����$���Qz�@�pŕRE3�Y�R��M�o��|�D�ж�y����f�Ȟ������`�ή2)cpа�퐜�Spg�w�����أ��&�V�3�>I��~
�l�`�?��&e���H-=����y���<��H�J�>���sb@��t9��Z���/!'�%$~����14�Sq����S�B���i{ݢ���]s��J��/О'Xq2Zߞŵ�/��I��B�4x"VM��+[�u��Y�^�9LU���=�|�E(��VjK5�K'��A�ݽ���gղÁ�Z���/mK2yt����I'��暼AG�1L��He7K8./�<�{&e���?dl��z�{��[��F��k�")F%��QL�Ǯ���24��=��OjB_���H�K�QfP'=^�򣨵�\�E��R��* ~t��v�w�d�@���6q�M���w]���2g2'&}AC�-@�zu�Y^+�^.�/�?�4�;���~�7�c<�P�,��F�K4�þ�k�ד]pfD�f�^@�ȷ�4�\uVA=������lRr�èL\�B��a�_��
�X��0�j8��a��&s���hQ�%����x@�����S��!���M�_F����VZc��5���<7��ԅ�uSu�w���Q���N4�ߗ��9=�4��Dq�����n�n
�q�����HCIY2�1O��tϐ����"3Dcr� e4Q�$P��L�� �>ǖ(�a@z�b�0��gT� ��R���Fo�-Pط�H�����cW&,�Hs���+Z �"/�c�&*XCt{O$���5��ڧ�Lb�ցZ_!�__������F�	^�Ug;�2��r��.����K�~;D���܆����g|��v"ȣ�B�*� [�\I��YP/�K�������M�-.a�!EjPq�gN����/3�#���z�G�o��>m�L��_�fV�K�ts*��S�pv2t������������|�y���v��UB�|�y;([�/	������䱁�<�F��ej�Ԑ������Oȴ�=�b=�7ճi0�hhq�֏�>Tn
����{���h��S��h	���@�	���l�T�a8�lm���k����Aړm���5���Ex�Eιh���BUx� ��#��^�)=���@�.�� ��AQ¥@����b�nnI;�1X'�IɁ#��$���E���d��#�A/��}ԟn4��a�r�B:��*�Ժn�Y�\��yҏ��v�M���'O��D 2֩%pۈG�
ղ�����
6������g��xõs:/T�L☥��-0ck��2DJ��N�����f�"9��!�Z��S����8��o���3�yb_[�4pFܼ��f�zZ2�;�޽�P��H;�T͑S�;�:QW6d�8	"�nT�kX袛-�A�	�&����Kp�8�NA^ ��r$�]�V���J���y��}a�.��tmR)��'z�z��:�G��e����\W&�� t����1+�|�ܣ�|��ww�=��_9V0X#w�]Ī�b�9��n	C��}��]�Q�*����1���%���EM��k��T 7��^��ͺ����x�vB0�"K���u�/�Nk��,D���n��5m5��X ��k��	��9k��2�?���2*I�kS��)
*�Kp�������^�-!e+K;;�t�hV��lP��Y�b=��=��dD�v�v�b�����<ȥ%Z:�G��\�z�%��=D����wYc���
�ɩR 43���	Ӟ1�Dm�P�3Q;#�01��"ֿ��sjt��r��;�}�:�~��re*��4��!��_�6�����`-JKXQʸ}�{��T>
=�<`�Z�	��@� ��	d�γ���:�%�����:�Sܜ��*ۮ�R��z�,C�����#�O�'D��G�[�$AC�Q�M��mY,�<e\����!�;w�+>��[�De�1��P=V�u�kC�<<?V��[��b �
����4����/Ӽ+*�:�]B@�h�{��^ 8���F`j9i��(NgIܡ��S�)�4k��-v?�,JZPk9�@+��T#��2j�ϲ�xF.S�A����*��M+��k�;�+Ëݱ������S���9d�U8a0�̭y̓Z���l������ ���(��qQ�> �a|��5��I��=�M
czz�XkS�C�ԋq(w�t����׳�Qc'������2�/�#�8`}���ÒX�	naEh�4ƴU_��{���_]��SyU c�<�C��m��S���CS=�g�S����F>��&���[�"���C/�.{*^EW�� d��\YoLi��O�h�� mخ��A�+X�� x[y�V��o������e �?Eŧ�_&s�ɪ�j�l����C\�u<yb�bv��c�a�(��Efr;��� �a9O?R��6Y�6:��W�%�:�����(�ذ�"*���~J�e�t���z�Ls�~�(���G��"@V�?cM뱚��������jp�'�����v!w��:7ǣ(�B�Ň�W��эΑ8�c�u�;�؜	_��j ��e�}�݆�:Q�!t���j��o��s�bmV�I��ܷU�`��]��<��� �r���DA���g�#���,� 9�
�\� Z+y!^G�aG�X�{�l	FN���s^PB��G���n9�zi �yg�(�|��T
�>5R����_�Vيs��p��C���\$/���*���f<B���j8���^;�!���Ry`2��P �G��H0��ȤT v��wj��qR�P��uՉ8�u���	R�vG���M�{�	�'T�-�j�:��Ƒ`�[e��%�^=崢�](�Or��C��@�Z�а;�E!��4��-hQ�Y|Hɡ��kT����Z"���m�$YCrK)���!V�
#�y��gĵ�ߜT�~2qii�v�7	�
�ߑ=&8j�M�7?]VK�*�D�{ha��֣�#�_�ȼ�t	؆��o4���]m�x�	7�ֶ����Rm����j�-�(j��Qmq��\?�.��m��@���V�04D��GԼ@�{ݣ�o�w��L�SڱῢY(��JQ�r��=�<�3H���3#������z<.�k�=���H���CՇɧ�ѕ�B,����e
kA�M�zѕ(�b�?��;NL �"�����B�0�e�(j��s8� ���b�~.��Ä��� ���d�e�� rQMxx����1{q�o�3�)���$��G�w����"��&���dr-s<6�� K$�C�����Kw��j�iN���4��Z�p�u��!&ZM5����X���YVLx|ddLyc�C���a�j�nFɖ�O��g��#T/����a/�u�u�1�3M�sl�\Կ(�xgj�r�:|�����{]u(��-]�(wa���:��	<����Zrw]e�O|_e��� 7�z�Xa�/<�ǖtV�p�G����&HP
V] �h��Ԑ$�CeP��6Pл�}c�e�i�;Nr�ki�4��$��'g��v��b���{v�۫0U=���o?����
l�)��mo	������������ĂC���v�nB1��*���r9�uW���IQj�Hjw�3� :�l�Q�??�/��[2+!&FI�=�<�W����5CZ���bJ#6m�����-d(�2&�$�!�:���_�^}@$'ey�m�Q}:>c�?�?��ԕ9���$x�Q��+��յt��A�Y���8�@�B2��v(\ڳ�a����PQϗu�g�� �h�f����2a������VٮW�*��ʏ���Ȭ�%G��Jp���r����lk[����y��Ir��~;�g�40P�O~�n�]��|i|�lӗن���X[=5�;o7�P'|[+�����|)LH�+�dȧ�c�;_����c���5�͇*��4%��
I,����PY��w��������L��O���v�,�E��)4�!w���ul�΍�30Wo3��]���Q!e��g��O�+������2��-�T6�ʎf.�n��9����#X�S pB���Q窐Ѡ܃Fӄq�p&́vjL�7�3lbAA;ی�j!Q��D��o5��h���Ws�TIC�o��)CE�{��`�������q~��`�ɩ�\�7���7:����'ie�ޤ�p9�i��ԍ3�BG�#^��5��� �I���b��wI�����ǉ�kӅ�d�#8�&*�ʃr�����M�u��k ��Ҍ�}�T����*��݄+�2�����E�Զ�I5�����oM�T�Gx�`�'`?2�&�]3���i8��Ҋ�I�4��� IW/4��eq����a��3��b�K
5x���j���&��Ή��nk*f�V��qFᡪ����:]�@�)S�J��GD�c�-4����(�Cw��`9�*�8@�!kZ��=/ފ�=ǾsEK������qUpƙ��|�{z&t��d����.r1S��^Y�i��ݠʈ-GGhGcf���J��yL�I1�)��%����F�<��x�U��܇���܉�W���l�3�����ű���ƾ�~�$����>�f�㚳R���k�Ȝ��ec�Ua�
bw��2O�a���D?�8�o��簸��g�`�g��i��=��j���d�d�~��r���r*.�`��~<��BN.��9�>J�mcǱ�x5>ƫM�m��d����X�{����SV��t�e^���h��br��q=�+'hi-^z�k1e�I�V�������!��~��X+�7��zF�� ��%HQ��I�|����1����+�y��h�N��K�\��`Ġ���~�h���F��z�O�Z�l�/��� H(B,5��UO��9u��T�L�k�.ٸЇ|:�!sj�c6�ح��P��*��}d�t\S��L���I�p'e����_��;>/���jE�h9�H��ن���Qo����s7 �?�J"6؛`��]K<��@�'��g)k���B�mJ���V�L��R;�xs���.
T;��O*��C�����H�+�d&�I4?)q���i�A�������#�]���Vu��v�ο�ɿ�4{7Oo]#�#��ⴽd�����p�Ln�J�����Uh+I�ګ'R̝��5?ő��+YsQ;�6��@ZQ5�r��x�K�S(�mSr"GF��o)���f~6=`f8d�����!U��<x_T^v�l�e58'W?B�o�;��e���X�F�І��Y.��8 wAx��xMO�i�6��ޅ?�7DҞ�Hy��&��0#���ݶ���ԟB�GQ��.�+h�vS�L�4��#:S���6~�@��ȏ��$��I�l=9�o�����>��p�W��;Ƀ1V>���\1�=2����dㅆ�Q�W�?&�ܻé�lz�i��ֱ�M�^v�%��]����(/����M7e2&#����A�C���+��F(V 7�C��+0g�Ĉ���zZ@��%"�6�r�UЏ\�X87�*{q4|��KU��#	�Z|.� fb`&���h�X�,
�"�b��9&)�)��ţ!�R����Q ��z3_�@�_�Y,$�(e��)�ۛT����C�v���Y���ݒ0�����$�,oN[�G`h=|�%hGb�V\� ĸrr*� ZHR�s4l�衼��2�Ŋ�S�a>)`Ly1N
���U�v��`��� ���p�ˢ~���E%���Iۯ��BCIri��C�VH{��A�k�f�{�,QF���Xy����Vԥ�+@�.������@!�T�TYҌ�o��t	þ$n 4#�MpD$2eI�M%q�����B�	�/����x*8Y%�֫<�rUO��B�4;��۹��w��F�	 wq���q�����C��j�����{e�1��{�����+D]�9a�0���י��l�N7,�W,�9�Q��[��-=A�7t��L�#�n���Ae��>�>�)|F����#Ȃ�f����a����_�)Ǭ�*ȥhmT"Dr'W���i4����dyq��H�mm��/'&༥:��>��c��{.
���/�@�%��*5Yg�R���엩��C�.i#�gp�1K{M��\��9~��w�$v>]���:V��2��T� Oݝ���;���Y��Y�4��1�y�5�~V�^C 0@��1M��$QV&�j�B��ҳ�2���n�Bq H�<�*��+�Ā��\wڢ�!߂%j���h$'h� �-��ƕ��[݂����S�����Awi�|73�	��D\\��m� ��3�H���ڧ(��%��Ƥ��8�m�c���x�q�SU��������}ӹ T�2)���e�y��V͊5o?.�q�9k�����J|��۔)�XBⴁ WyLb?�>(��A���Q;�2x��ȼCO>�r��_��/�%E=+��8-��.��ĕ{1�rsR��d���|U�����ad>D83<�$n���Q�Z~\�@4a�˙'�I�*����%�*�:��N�(���M��ه�n������2�h��9�7�A���M���4Ku��T^(�m������Elr]��<~&�Ix�p7$W���sP��S��S�ײ
~qJ�=`��Qa�-��>&����*K��P��K������z`\�L*��rZr9�1�7�r�1'��弖�H�L��l�dݻ̮V֥-�M�7\LX���p�i�#S�`����}�bD��(,�f�P�R�7gw~�IO�Ѥ$�6�T��Nt���nkS���/���#u������f�E������dug�S������%�x*���!��z&��a�'H��P������q>�kp��t�\�T�sߧ�Q�%���j�&;���D���Z%ݥ������b�cl�8�s8��ǣw��p��\�v����@�ݣH?w��V���g����#�|��Q.H{
���'�!�a!����;�Y��\�P�s�:����!Z��[p�j��X29kMW�ç`m����oqtI{G_ED^q����
����f����6pzr]!�hoֹ����?,)�ͦIz絗3.q�I����Q?�k�\�8 �;�4g�DL���`@MԤ���aӢ��J��	�V�^M�aNj�^}=���aƼ���ShՏk"���NB�4P&�R@���#��v1�Y y!�:��
qx���
w��'B�1�u���29�	�W MC�-]}��iy5�3�� La�J�ϔ�:)H\�6Ġď>R���=d�u�3M:�[�(/��Y�����Uy|��S����汝OT�e�����G�g����~��!ou�uy-)	�Ҙ0�X���L���国<\�c�����5oV/Y+S!���@ܦ��*c�oQ�/���Ws�:�t�9�n0푯��(��i.9�C<~m��Fi�ʖl�O��0��8t��'A���ۻ^������>�؃�S���QVE �X��~��	{��AmV�9R�:�;Jm�Xm�3���L��4��g����!ц�b�(-��2HpTa�6/ҼW��4J����P�H��<"�)(��G�����ՠm��-<<�$7��8�=���!�p]kx�N���m�1
����uK���a8�o���d\����L~V��s8Q���_U8w���r��3�K��5�x��$�4e	7���o��4m��b�z�@Y6��v���� bNN[r²L�O�_����d<�ėW�d��h��yOA����V�+K^:�:ݝkR7�d��y�l��?ƚ6��!@��
KsB	b\�Bw��;N��� �N�$8�5F������D�t�J�k~Ou��C��R�JIb��A��� #!����+�J� ����mO X�]0�3�C�I�d���ga�_�ص��PH�oq����K�d�t���dlѡ!r%�̕c�8�y�՚S�h">({R���UxxJ>���i��m7���� ��_���qI�>���S�y2h� ����'�ŻKl�h�j?�9lm��Ӱ�m���Ά��#ϰ3t���+Di���~6�{>�X=�,@vWL���l5�� S���o�[x#��Ik(�ㆦ�t7x:!��8�����P��pe�<���n��l;�����lho��������)E�f:�&S2��Ԏ]TQ�[p0=a��:����,S��UU�l���05I��P��&�F)���JԮ��妐�9U٬��8LW�2�I�����j�+���a��1�-)ͻ#H{�ː�G�&�J��k�  }	�� �����ֻ�nF��f��~p C�&.GL�&�a�8w��z�߿72,=��V+߽�I��:rU��R��u�g[��q3y]�v��4cN4�k�&�Q:����j��CP���9Q�G��u,�c��qB[���n�-����+���nh$c\^8-S�x�iN$!NQ<�J��]� |>{2�ZAy���_:C�'*y7Kw�g��5qs']6%�%c�vRA���❉V���Z|�/4k֟��% �E̠�F�����O�/�"�2"z1�"�e��v�����M�S.'P��M�
(�i�1�\� ���z�i6�5�gs��D��x�Z��Ŵ{Z^c"��u�Nű��{�s���P��qV�)���(�JuǱ�z��M|{Xu<��_B�}�/k$�$Va(���:���w�r��Z�� Q�se�lhx���i{ώ,k����z�y��SQ��,�9�)7\>��=�R�Q�R5�@�Z��xg�U���s9p�i�u�¼ںV�~���`������lDuG��.l����V�wd�	������������6�WK:0��N �nʱk����ߵw�՝��u�O9�-��_�}��}xp�CC��Ք��M�E@�3�a%��0|��u�/�=#��q�C#�s��g��(r�GR�@�=�&׷��~��~�� �h�)L���HF�
Ǹ{�%������c� hh���}�Bk���aA��U�Czm���oX�4>���g��bY3����,�~拟�@���+�%��*.�̛t�5v}�E�]\��P�l�-����ˁڣx�RЗ�2~\P�=w��Lӕ-���)n�E�}�����J��7���W`���ϻ�\���C���߈��D��'5�����~���^�9@��g*{�@�(��搀1>lK*�{$\���}#��v���Ε�IU�I�cz��M�ƬzuzD/#C�*�>�=���nP#��gB��J7������o��f<p��Ì���^��zʌ�P/�88lE������K�]��t�|��\��k��	l%�V�gQ�����W�� �0>E��wǏ	(/���`I!��&Mf���(��1Nk���C ��ͿV�������Х�#���} �*%8��M��(:������u�m���?��j�MD�ƈ�-˱X��s|�:�����m/� F5�cP�-��ro�i*QTBMa:Za�(ϬF���7�V:�p	�1�A���%Pb���x2̟$�]G�� ��
١⦁���􄆯�E������c������o�j*���b����:*�X��T��k�i�5[(�q�uB~4v1����͠�7�[�B�2��6�|+����Ǘ���1���m&
�cf2�,c���GӤ��*�@�x����rnrO�T\�e��&���O}�=?�%w�l;B�U��yz�هn[Μyi�xo6ġn����W�ȻY)��;� )�No��g�=�yd�mq�.9����O�ǋ��5��o,�嬛���
���"�\}Q�U�կ>Ι�<�,���Ch�Ċx�m���6k���P����I\�Ij�Ow�H��w��=B��p����J���qY��( _M���)ˑ��o��QFt����b�"ד�UZ����h�`M\<��x����"�ң*����I��cXL����ނ3G7\�>�&�4H�0p�*�)ɡ3a�h�g��[��g�(#���SE����9n��]z/;a����k>�q�o�7*0 ���@���#ǉQ�K�\Eh"��uc.+ژ�MT�8�Nف5�Z�o�u���O�I���M�Y���D/�cA������`�Nkq����HV�xS]%�n�����޿��}?~��o͕�` �ITcz��9���.��.�Dg��%\���qg���=�H�n�]FÊ�;���o��S���6�g���fa~�?�D�(Ky�¢�h�7D��"Y�b}��k��X���@!�xS��z^�Qg�&@�#����u�у�� ����$_��V�  LUܞ&'��e9^5��C��#.o`D%
��i�
�����S�77��ybZ��0�#ްYǹ=�&f�=��	��T�7e1�߸Y�f�@�v���js�ޜAq���P���<b���:'f���-����8�Ax�⮵�V�ת!��}�{a�
:��A^qcr�1B����#�+]��<���<8�����Wxy��U�1>��w��8�IQ󛩏������c1&�ɦv������M��a�o`�V��oB��by}��x�����NݙD��-�Yǉ*��!3�
,�Zu��`�z��~��!��;p�r� U4�~D���!�,1L��#�afS)o���L��NM�8ję7^���2
�$Y���PF��d�	{�S̶ŝ#n<J�qL����j��U<�:՛�J(�P�΅1�Q������EI����P(ИO&���x�Ú?@��DX_͢5]*��c΃g�1O�����a�����G$�Y\�;5N�����`��B.4`��D�롃����L�V�/�� �`kc�Z���U|t��=˰���a_�f=����ɂ	�n��{�z�x�X촷��u?�g��b��j��#te�b� ���u�Z͵{�0��N�{��,��^��Zwb�i�)X+��F�^��[���p[.��z�t��5�r�d�f˦N�|����l�ǥ!{Z5t8íI��Fڽ�@.�0���z;B�u~7��h)~���1��o�]L�>V}�Z��vP7-���RIGhu=��n��,��0��[F��iT<�#���2����Y�{Z���\�K�����l�]݁t��U/����6m�����]����{�Sx����;)�v�3��ڴ^�%�ۖ�@P^OV4pz�A��'C�R�vݖ(*#֟0��Wcj��K�Q}Q��J����F��jl�BTȄ�M�i�%�XM2ԕ�L=��e	�ׂ��;�+5�]�Z^�C�J	��a��%�`���nE�g��&'ܸ�'p�w��x��&����avVa5+\e]�1�ؒr�D\<.H4�K�ꝿ�{��Z������.%�PHű�e��ш�d�#ːҍ�v
�7#�5G���u����&���=َ��g�B��^&<eo`f���.���m&O���T�o"��%�Lʗ�]��s�,�SV�?ێ��.�=�r��A�gӈǿ��-�|�r;���ᵖ.�t�*{���j��rNЄ�&�X�78v>�?���)��X����m2J�C���	��>uI������pNϪ�0)��7�1�������#���xb��h�<����%2�7���s�����p��E��=uOl����У����6G��۰��0���$G�7"��:�+4��6��[(8������͝�a�%?jλTp��t�����-B3�2[�4�^朌V�5��gD��\(�K7Vs������cXƂ��O�4�fq���8$�o�r�� 7��M�c��]�.����#������Y�L��mE��q{i\~���ߊ�s]@��^�4~�uԖ���A���;� �o@ވ�ˀW�up�)��y ��1�����1(��B���3�O�������ئ1�]f[���y7�0=k���O"P�ڟ���i9��0"J��/ҙ��39���C�u�4S���;��^�4/-�F�i�'����HLb}�E��ث��^��;��W�J��x�)bq��
�b�ЧUˠ�;FZ29�s�y��&;��w0P��봹v�d�1\�&�bĳ��A�`�2ҳHd����C�?�Co@s)�g�]��V��d^���p@A��co�����s0�Q+���:���5$�N��M�Quj�Q���J<�5�P���e�
�_��4�l,/|��g2%�w]�QS�!���n�:���Z)����LX_
<���yE�( yD
@�.�W��(�������G��NGm��RB����Q<�Rh�a��5��Tۋw�`m� >V�[��؍+�:]'�qd�nh�E�k `�q���K}�c�Vc��s��I�?;�V�3}"g�\���ޅ��.|C �):l5�lp�^ƴ[��0{ޠy�:����KR_�b� Xd�jw�8oŦ��V[�ŝI򘂕�����Tt\(F����潒��Ө�Exq\�V#jy�^���wa�*5,DT�]4��;�[�E0�� 9�*^(����J,�����b@�t�u�8��ϸ��E%vGҁ�Z�g�̞v���V ���I�8�����Y�� ҫU`"ц�9�g�iP��k��a�
�"B&���X�Ⱦ�vS���ܸ���)�~_X�g����m�E��3����J	��n�n�X�'�Zs�"7tT���������\�s����{r۫t4���TT���Tu`/���9��.V�?�S�����1ypoE`����!݈\+��Mo��$?��-�<����J���i;ӝ@'���?H�Q��I�W��A���?��� �IemZ{\����S��٫�p,K�ÿk0؀e\:�l�l�1c&�&�G�Aw�H�|?4�3����a��GF4�ҩ+�b}�=BX̥�L� m�,�q������h��f��:t8��[h�m�WL<�zZ��.I�odQ�a�E�^���04��L��Ǩ$��{nl!dgI��,���,k��.�|�U7�l�`�(%p~-�m8����͇5�K�Q��Q;��GM�������?����-q4�7i�u��M5LmH$q=b�%6H�D
o9�{KM.b�
�V@EXm�sTO��8�޹��=��q�ed#� 8�ÛC��`�Yp ���B���?S����On�/~:��X��k�\��Yzp/dj�):*��!+�8;Á�QȞ�Yx8��w���%�.�nE��ed�$�����Oz���ݎ�f��"m�yW�S�S�~��+�˱rn���4�k����M�f�O
�T.�̩�M�4)3A��0'�^"��������b��n��C����{$�������ں0	j{N v�eRѤY�����p�E�Kh�`r�	Բ��>ed#W��$�ɎH�aKA^��	��c"*��])���/a���b��E�<.�o`��`�����LCi̠κ��p�k?�2��GT�/�Ƹ�]�D�L����B}_iLiE/�����HN�Nl�s��.bGOO�aΦ�1��n�n�f�&̺|tJn� �D_ʖ\�w0Бn=�α׫cUմ�z��� bsqx����~Z_�~F����g�Ƌ�N�����-VS�O~�⎇w3�F��_T���$@���B`=۝:	�m��.n)��oؒ��@=�~o��v<K*���[Z�'�tLΧ3��c���l�{��_e�����DaXO.��;�����n�Rr#��A��.T=�k�N�MLkKfa�t�=�zNjP7,�E��|:�^}�@�+v���Mh�X�#"\	���Z�>�K��S
t�]���8!s����a$k�d�9�{��0[G�{[���=���A�c�X�J��"�T���7C����$@�X�d~_�t�%Gzs鶺^h����I��	`��r�s���@<��s`���mo�Q=:���+8:��K�&����Es�%��<:;G��Jt���$mIe��*T���nk����I;;:�)�M�����a7���?�{<90��?���� &��I� ���O�a��������w��fm�#c2�˜�4�_$+ʨ�h��D���⴯��V�N�&^Ł<��	 �:���@���e�dU�/s�{�-��ĚS���2lyB�2o��O�2��t}�)����F�/*�8��d��
��`q����u�y�ণ�C�hJ�U/�_���M�sB��M�������2���7 !�>eaDps"�\$�o?��$Q+OO�6���$�J�;$.��Q}�~;�p`�
'�,uhY7�h�L"�p�3�ׂ���Wm��)��M�L��bS�t���D�*���`wn�%:���x��A��Tt�'.o��+ω�B�� �$@�6'.��g��\S�f#��$������۷�ڳґ��"$��kV�bgb���p���ЃpDL���7���E#N	��13з�9��\�sl����0i�C�	7h�.F쇃ۮ��E������z�S��>��|a��NOCyJ��i��ː�;¦B�G=ë���q�k��b��YM�U-��<����<Npq9��9>��7���~4ƣ\7����kK���z��e�>��-!��S�áw '�Y
��k�J[RũT.�a�>��%�Ԗ-�����l�H���X��5�&2�h���mi��S�(��B#�����"z{��ܷҶ�#���$	K�4�����I`?�>�N�ky�vy�|�:INàR��J]����PW�^Y%>V.6���06Ã�,���#|Ǒ.M��J"e��ͨ�_?G*pa����g=�PB��J�p��OF\v��;�Gf%'�J@?M(��<��~�n����v&�,��!o���u�eݑ\W�Цt�Ȅ/'~F�_`����y �� �n�V�	����.4:/T���[U�0\���9U��J�!�Sjr�u��K�m�f�C�l�CK�4i��Ϛ�uΣ9-&����FA��������ZzR�a��R�O���o^��qcB�@����H��]|�p���~c�.�
U���'>�6��+����s��g��1�����X;.��;��5�kH0�w���_��>��A!�!�Ӟ��I���Uz23�r8�@�ċ��X���ٱM�B�wI-��a��KG�Y:�HB�}�%t,�>_�-���xa(NsJ􇆴q���=m�-��@	ԭ[�ed���j�_�\6���i��I�+�����k��+z�3�e5�Yx������r�(E#�մg���.�<wm�x� �t
RM䮕~�⋵�À&7���ā�M�)�(�*�ݢ�����O �P�A�N���b�}E!��Ni��p�%'2+$�Sm��. �^/*�x�u��{���$t�pH����ȗ���nK��L�!o}���u�9���on$� ���^����*��t����H�0�Dn4�e�)�F��S�*��"6�>�^�&���n�R�1%��w!o� 	v! ��֦�Cs��&ɒs]� PƼ`r ;����ޓk�����+���O,�$����wz4�>��۸zn�4b�������Ϳ{����}ޡq-o�z��ab�7u�[��zWW�'K��͞i��gN���wU��$flgxө� ������g�|�7Ϲ��%���BXY
�Bp��i��d�'�]>�#�_.��87:t?.׵K����0�:�F9N�9ؖ�S��%��L�T��Ew��O��ں��� z�>��;0�_܍X��OeW��|-8Xk����������_�X�-#w�� �O�=�bD�kD���7K��Jn����H�w!!���G��W�j��L���L'�E *uG᧸	����KͭQ��3�e�{�%u���G�݃�W�;�OYGD��N����Ќ|�4�-&ZX��p�|2_��R	y�>�Va�~���᭄U���8�������"0���ǻ`NT#�I|{�Ъg�蜜�i>�Z|E���OY�����I��� 2����-_�M�K���KQ�����̓������AiJ��v����^ �S��ә���m���ݺj��Q�~�;Sm�߳��������&�|�ųf
v �F�
/�~E�aP�ܝ�|�y���?����f�+�`��#C��1��7�Q���%�6������,ͯ�a�ct�ѓ�� ̒艢
�؀%�^q~�GcN3,n��SR�	����oW���eՒ�^���q�^b��U�o^/]����|O�/�젖�L�5eR�!E4�؂�<0��� ���Ն�J�/���Mb���њB��)x`~�S}���鵏g��d�{�h����M������OoH��KP�r�j��k�/S$ˉ��웯ZџI� ���	��x��������΀����X3�ˉ�HƮ��v?��iB���'��(^��C1y������eT�,���5�fx��c�wIVcdxK^0�y��h�s(��o�W7;��xm-ڼ��GTP��oH"V0
�l��y��0~�T���v���c�	8u��@��H^��L9-2��ߓ"���)H�ȧ�jQ�i�?SLԇ�"�F�i3�i��NW)~�;���P����//~#������q�&rX���>e؋��o+^/��AC;�%ȳ��V���I�����$��������'W�/ݵ�Rg��ِfh��Y���ܿ�I��Y�UE�)��SZi}�����V�,����=0����+�~Og?VoۉυC��X��q��a�Dǖ��-�7�GI�磡qLu����N|?��#��Bp5��B��4r�����w�^G}AէMgk�1�Oƕh���O�O3X��Xl`���8��;��ȝ�4���r�__�v��#���.��t�*��~�T
L��K��/�U:֙#K$���R ��m3�8e�����t�W+2�#� ���F�^��۽b�gB*� ��9ߑ�Ս�T�Vш>Q:�ꖋ�b�Na�7���ǤX".r��z�K�J�Q��jFQF�*;�����N\WO8�W����o�����P��eH��h�Z��g*\C(��۝5ån�yw.\�G��2}��ڤ&���0El��5;n���,�¾L���H�_���ɖ�D�G�#��tk�����j\ n)uN-�Mӹ��4A��U3�Fg�G��M���E�-�7�&׿=t��ܓ� Tuff�[��´4���D�v�Cp|zCZ��s�b.��r�=ǊX�lM�t�`\Wȸ�c�xo�v����I��#�|'I�<��"V��4�)n&S�m���cʃ�e~�"AB2��v"y��`�ai%skٻ9��}�+�bC.�F2,�<Iv����ߏ_!NTi��, �ym]$.����>n6w�h������\ q�A��=nn4S�����g))�^]so��5���.O@ߡ�,�8�F9W����������b
1	��-	�ЛT�D�^�����I����+h�#��q���΂�/�54�~���zh��g�v�]�uD�u��t$������,��7K-H_Ha��XRV��f�⌧l��I��W
,ݎ��`=�BT����A�������������E+F�J�Ne�A�[4�q��gV�R)G��}� 3`+�� XaL�h!�B��>�v�[����E]>�|N	�!��1J������S&�#rH�D�F�ja��k7���f�'*Яu�N��-}�4��[d�<A�GL����;=M}3z�`�T=w֤Zmm46ё���CA9���^��&mc�����v�e5���sT'N��U[m�52�{�h2ac���c#��V���<�w�T.��|��`*����N��FZ�	]T|gX/�����T�J(� ���٘J�CE; =���Y�uyk�����p�H��4}A1���X��o�h���G�����A;*��.���t�o;���Y�08{���"��'(`q,k,����Vg�J-�Ir+��q�Q��?�ڸ�:���HD�o]�r����x9>"�V >���������	Ы	�Uؽ��He��ɢ_7�#���J�N4(��f�]E3�6��#��-� Is�JȖ-_�,S��Ц��WD~d�X�g��L6P�iR�����e;:Z��;n��%���d(;��.4��[�s�s�2�º�O�� k:]8�9+��u����o����ީ��ԅ�K���Ke+ߪ��躞VKa��L�)���{�U�8�r��1�N �:�j^�Յ�]ԟ�����.G�Kʳs�
����X:�����L�Y�	,��w�*��Z� �?�M��u}�cwv�l�Y�T�k��2re��
�`���ci����շ�Ě872�v_�xH�'��cg�@��~H��r򆂵�-�RtE{M�� ^F�����f{�d���ܯv�
�R�)�E���w�rC��f�#��[��Ҽ#�T'��zM�Ig�0(��u����*&��pQ�>6���[�����w=h�rL)�:�V:d����3����\ �m������g*L�����iH�a��m�Αm��V&|��Ă����6m�x2��>��p~&��5Ɇ��Ƀ<?|��u�_Y�Ĝv�Ҽ�A�ހ�Be����V
�s��`�R����fĒ8�KI�Y ��1L�9����MUXO��x�1?�X�b�!G���� خ����j������� :�F}��i-��%�+��(��u>}��Ȁ[߯g(=��vh'����M��k�6#���An��^tg���'NX�u^�\N�Z��l�/I�K��1o��*o�#��t?9���Q�ZA��}��g?�;�e��L1΢� �K����F�@�E}�陆(N=��
,60��[�޲DA������]�8�C�Ӈ0K�dIG���n�V���`���}��@��C?�n�27ZHO��:��C��ϛ9���ͺ;�9�Q=���ru� -}Q�1UC�	�t��p*�3�~(��wDa	Ս	�@Q���ٱ�����+�b�-�'Z�ҌZ#��q
)�M������X�y�o����8Q�^%����3߻�W��R&��d2u���K)>���bA� 
+S�zOROv�+xZR���IB��N�� a�]��&j>fB^����f)��v�"���-�vo�;�N�H>��DX+6�Ib7��+���>0��9�g�#�ڹ�8�o����c������H��E�䇃��u<#�)o�ZD� ^T��L���K�V(Y,Q��V��@�H��Fes� �����1C�Y��*�Oe�b|�a�kL����u$�bVp	ē����fvW�Yu!߲P�z���3Y�>܎.B#~��S�͟�׫�H�E�c}��m���ߪ�\��p���X���QFtZ.������-�7E��0����I���HYN��M�%��jA$4�0{1~������W�����x�0$���Cm4�S��")�D|�N�m����˓��>��w-�Ҩ������E�S���r��)�^�D4ǅJ��7�1��O8�Q~�:$�o�2̨�����CDۍ"���.�3Xiyvu��pt�oH|���[ɹ�cfj[cf=ȶ�Q�ĤRY���W]�WmcԺ+�A{��D>Ŗ����h�f����B�HV��X�U*{� t:�����l�������}e!�I�Ä�6��0G �f`5��g��~Аl#��g"@K��ZG��p �t�E��}c�X7�^ ��!'�d�����aP�w�;�������*���o92E��NhoDb��D)Z(��������ը���Y���_�ҿMw=�N2L½LA|�k�4Ӭ<�3�!��D�PU5���j��&�$�S�l�u�h>�%Z�	5�ĤaP{E���sɩ�|-�){�8*�M��$C�p��3�Z/�$z&=ߥ�"�d�9>���Y(b7��oAl|�#G"\�� �Um��}�O�/�������N;�4w�h��lW��	�<M<�3��
oFBE�*i�@i�{7ox���4έx[� '�X���{��V��	�fVA�ɇ+I�Xr�ȥ>������Ș;�F�%�h��T�9H�
�J�2�#7�	�h��ohu@0�N\��KhgK�aA�x1b�J8�G<�Jd*;���>nX������#�d������b��ғ��)�Y�!�G8�w��k�Sޫ�.�\�L,��&
%�OT�;�^�B-����̎�8;��8�>!�8z^nS�ik0h�`E��P[��3�?�y`k�Q �?�鐗��0�߳HQk)J�5z�\�#���kN}q0�r҉�G���3Ĵ6�I�ZN������g�H�g�G܊�S�V�ڠiÀ�XA��	�w����]!o5.pK���U�F��o;+�1?���!���� NyY��L��3Z2�+]��Ђ�/�� -u���d,��7�m�)6�!?�D��&���A�u��)&	�F�O�X�F��A��/4�/Jh���6�&��ںY�6,M�/�K�G���=�(t�-x�?�U�𾋚�Կ�o�Ϧoy��Sqr!ˀ�������{C�1ƜR� 6��-n�Ve����H��c��:�pl�Ko����+�aj���T�Qa�5?;�G�1�mG�OZ�OZ�Z��o��`/���z�sO<�ԫ�(��3G܈C��Ɵ��/��L:u�xt4h�i��Mf2-�p5��Ql�����y��kD[��u٫c�k�s_��ۘ��i�9�ٛyj��E�����
����Y:�1���:�F�)zQ+�B��1;�?���|�%9�ꒆD�#��P�A���X������ET���O���ڙ��E�flx�wS��O7��k��u�v,h�u�f��Pj]�V��e�e�X#��$v�HP�Vv�k9�yj $������0�� �D_u�/��+gn�0��*m�$E}@�=�$�"C���:�d�F� 9udH��6>�j�{G����3��x���vU��q�cA�p��_��><r՚�skA%Mg&��8����w("{�Ԃ8��J1wd��N��,�h��ؖ���J}u!���> �7oI킱vk;$������h,����/��8��w�N����Azކ����rC�6��z����Gn�� �s5�Q��5�H;Q�V8�H���!n���f��"�D������.�C>�w�>_�{@���Ρtj,���M��(�x�4ru_��+ȩ�sJY8iy��$�4�w�uy�����֫3 mi�j6���P��r�����ĳ���>T�jUC?x[�Q��	�.i̘^�3��ȥ��u�,V6{Q�e�)��q�0v\P]#l@�&��,��3���7�<�`�Q�%6���QZ�@m�����|�q~�1�\�3'��&���͐&�G�S_,-���q�
��?ⷥ��K$4��ЇW��L�T����ء���n8� 1&w�ؘ�j�7BGUk�]��.Z	��O|�]��W.�xG̯0�l�z�ۈ)��g���0��
�E�ej�Ǘ�e�E�j�YK⢔ࠢ0��;~��C%V���O���!�P\}'9|i=s}ȷ(���C�w�[;�E�=�H�ZXcK�+�(�w�
����U��2��!�5���'��h,٣F:�����j�>��� ����6� �N�)��7� �:��ȍ�x�����Db<��Ǣ!�̿qFє��D���%���4L=�w�.h��89#���M!^�>i�Mz'ŝ�s��x�W�=
��o���R������}#���4O��D�U���J��J,�L�	�潎�ůݿ�U�s 3��X��|dgjp�:( �\�^�ym�A�S��u�\ �
zJq3nh0�@�$v�ܔ&'��G�x1!㟬:CT�Ԇ�Yr��~���#l�6�+p�h�����.��+JA��a��W7#��Ȝ��.����T:}�ސ<�������oF����q�IC�)0���nq��5,�x����P��}� ?��i��AT�/mmp6���ſ~���֙��mܾ���w�hD��	���W�\��~��I�,�u���]�S�/�";�M8xx�O��;kU�NT�W�W��4�?�F�V���� �IZN�*�b��������ʡ���J#�k)�˖��ɧ\����+ע��&\��DWJ�����=@�F[fab�_�
�)�-eT6���̇m����C���ғEI�ҟ�G%����t��+?�(��@ӑh��$b�/(\"��K 6��R�u#�y���\�Đ�y&$+x����E-R"����g]��x�]� _��0�*�� �Z���ԋ� �1�̷�'��g��$j�(6����/�s|�Tm4��z���f{W���	��Z��_#�G�j��*V)��3�3C�?�?�����A��W�>2� ��Ok`q���ެ��5�!Z#>�~�6�P^6.fCG��Q��uS� uxL&gb���m)j�U�Ǒ�@b���{q�g�$D\����St M�$+$yH�h�ݟ��#0��2��ø�y�uC�([]�c��}�!�-�ޟ�]�L�?'弬wh���7g�3<}�.Nt��7|�sEԥ��na��@s��A0X��KQ�|	J9+Dʆ�7}
�./�*g��u��p,[� �8�UYE���x�H��T�qg�a8�%B�t���z ��A��d37bG���st�9u���S�v]E������s+�''&�7��\D7�]A�:-܋��q����!�n9�k��Ə�iѧ�JU˓d����=��W�bZ��{��11 :�vY������c �����iE�u�f'`��_�$�X�8+�V��*��X�g(�H����^�D�_qLX�v$w�ֵ6��C�պ�F�_�5���T8HxK�f�#Jâ��gye�;s���N�Jx���ʞ�J�خL��C�.����I~��!�5����쐾u�C�Q���b,W�]&e���9��� ��`H�Sz�VcU�lC�b� r'I�<��f^75p4P��1YTa�-�e���� K��߂��DDBs{�#V��p+�,[�j�;�Lw�%�`t�Ӑ��`gӝR�P��H�LD�bk�c������ٽ���oo�]xk�sޡ0�e��f*���V�>���h�c6��v�^#а6rɇg��[ޕyL��ӄ�S#W�2ؿ��K*��XNݠ���D��Y�F����T����(W���\��2�6ci<�ES����B��‶�GT�u�(;̈��t�)4ɶ���H2|���OE�w���u.�dב��m�0��7&F�L7J��Ňb�}�`4��X���bE�I�D�9u�ɪO�v�9Ż�2�f}�a�t6+F�|�h%� ȩ�0�RY�nv��T�)�b<����3K�ݢS�5zĪ���!a�6X�:@��!C9]��,�V�M���#3�	��eM������u���<4��j3��Px�0. �A�N��J��_�f���Il���
+w(I���p#��������%Ķ`�����
`����ï����G��h���֓V�^�.I��f b���p���N���7��|�jft�J֋MV��4�iŪ�mc���J���Q��Fᜏ����X!F���'��I�W��Q����/�Z��z�7GU5C�%i�Bᙫ���>/ctW����
���y��
�X���{i2�a��"�X��*����>����*R��y�*,�K�/KkgZ.
���9f�a@��|z��oȡ'����P,6�l
+H �Q�����W-v%��H	����I�=��i#��l6������?S/�ix��N�
*��ެv+����VyQ�5F�T���b┑�/ax.]�Q��0�����[�.M+�'0V}@o]�`�޷J�	R�I�32�5�\�"M!E���fߝ��=�:�1���ר}�뚪������{uP���2N��#9rn�G�����R�hC|�M��[��a�"0b	�*Ξ�^4�(`',ʚ�f���W�d�2�*���c��DB^^a����Q�B��Uh��C�D��k_s;TA��Jp�T0��
O2Q���� �h����c��E�(�t^�J\���k5�c�����ss�>Ws�����ǲO���gPkDq)q�{��E�ߪ8�tM٘�$� ѭ�pD-���q�Kf���c�8��!�[L�R3֕�o����;m��H��'������8҂v�I���9"F�z��G���M�֝^~a8���ek��(v��L͌@��y1Y�١q�hjcf��^�J��+�Ԩ7g��Mi�����'n�{4k��X�/�d K���A�̠��v�ߜ����Ew����{xj���*3V.Y`.���ڔ����%���',�bJ�Po֖o�gʨ叐�y[�'�_;ui�.f�jX�e�"�d�Ȇ<�As+N_)��dw+��:1��Y��hW�\$���/�u�^�E`ڮ��hlMI1��j��&m��˥�P]�����TTdZ�����ZC��hJ/ˉw��k ��I�����mv�)E�)�  M�����]��6�D�E2�}r0 ���K��55977������R�'�|�:�<�y��~�e�y��sk�(��N�b�'l0C��f����e��q����>��`��#�*�HQ�)�;�VU��~M"��O�X<����U�����J����>���R,�o����ݓ�o>��T��w��w���%`����{��\)L�/Zr�k���Y�ff���{_ ���`)kLb�S�D#��nV������m����F�{M�v-7D��IL���y%�T�HS<��P@�$wQgb�������K���nِ�fM[�t�NL6�h�֬_�鴲�V�,=oL	w�6f�������Hv6�&���'b��A*a�W{�W��>	B�S����B����"�k	�P㾺��31���߷�$h���p6!X$�|�qA�<'�g���G]Q�Ӯ���m��I��qAtd)[i���� �@f�dJ�HC[T���ֲ�o惕��q��Lz�`R.cm�Sb��=�)ۚ��\�-���E��c�>w��`�+0�TQ�Z���wx!�ٵ0�M+�������_�JL�Q�B�70�-� ��sJ��q��+&w�,Q�ӧ�f�r�T�en[ۥ�����9����]�T��~?m)�4��ᤀ�����.�r���u��l[�+�h�iU���[	�KV��-Qo4��I��Z�c�ȓ�c�&�KV"�Uk�i��ѭڜ���%U��s��<�^�c�:O�Ͱm�����@2����Ѱsv��-�V���-���n"ԟ�H��� �j�w�v�7O�*�)M�Cbds�}qoN�۶�]�d�t����@9�ڊ��{�6	 ����������g0�@�[XK`�H�6��M}�(Pf�œ[�O�G籋����cp'�c��b�/,g�'�%cw#|��*%�N���Y"Nu�D��Fʲ�\�;k�)F_��)�o-b�;
0�}o��8�����*v�ן���N��I}"���s���
c�lU�ut�'�W���ۓ&v}���eg=� ��H�گ�(Tx���Y���� 5@�S(`7f·�L�Ge��,xo���'�B -Pt��1y����og�L�]9�tr4��h�ɜ��i�����R��U���2�\8�Ŭ+w!�%� ��^KJ��R��oxUӠ|�A�u��9H2�lSNW����5��_ޓ�y��� [��־;˞����8�Y^?���П}���ˑ�[}s�Z>�%�*��2���������^̴�l�eSǞʩP����g=đ�Xu��������y��섽�ͽrd"A�,5,[�{�
�	�ش�����R(g���f���m��>e���sT���/���k���WO�H�(�Ph�Rg���ޤ��_�\�K�f�e.k�}q~U$:S���RPxMG�7Q4(���_��;��T�	3?Iuc���é��Bt���c�xp��a䍦yj�cF�����N]���{`c*ee,�&"C#s#@�e?}�va��sD��h�D�6�8��I���]���@�5�!#��D�c�A�oR���o�f!k�T$�*�m��&T��%��,���}�="�)+d%�t�6��MҪ�{V���W������*W�*���4o1Ƴ�j�
7�-j�#ń�H��cW*�UY4
NX���ΒR�-��z�P�)r��Y���BF[�txM���kn� ��@�����+*���2z<�嘮3<󀌖6�@E=��<�D�[Y��g)?7؋�f��kk�?82�㓊��l�6�\��ERI��m���G�sP��[�p����1���n�p����g����!�h�0)���䬼��v{i����bJWy	S8��QG��߅����g���#���D`ܿa��ǋyi/z�L�(�b�!�CS�o�^�f �T���'�(�~	����5g�2EEs���G�î���TV��ma���]5����D������9���j�]�؉�F�R�SBk]S\�׋���*�|��G�I�'gD�V�SC:�U����ڏ�s���َ8^N��<(=@	��Q�=JL�EN��� ����$�K谩��Q�,<\��ߧ��W���
>�3 ���W�w�E^]T�J��2��fчr�����EDykď��CRr��і����̜����w�J;�h Sܸ����3���'��J���Z��!�R2��*�}'|ur{/���Hp1� m��6�m>*;Z4�x�Z� ��R���T�!؂��}�/�����p>�����VFg��L������x���3�eM]������%e5�Bu/,���(�В�w�b�>������
n�G�7UG�����8>�u{��͗w����!L71�i��x�h�aϮ/Eq@R������L�6*�}~!��s�L{�_� �����ýlC�2�$�]��ݪ,����8���1�QA]X�˅���_��Q�7�u����B���?�Ҧ��Kk���X��?r���(a̝Tj
���墫�(��I��O��P����\':����ML����H����M�B/}�G��]f7%�H�MW���R�6ߒ�&GOzm�M�Z4=]@��]��[0�����j���^E���%C����>A/��0Ԫ" dtHv� ��Zm#^�n��j�͌'�6�������de�Z��8��&U��p�?L�4G�qE=�����0��ը@��"t+���8���v�($��e���o6ܽ�+� ص% %i�i?���3�'�e\�ز�8JH9툐T�67�x��惽`(0X����jl���g����#/ل67�i�G$�w5�2wYw}U7������ޡ���g���K1vZ�����u�z6H{	{qw��Z�[N1�R��e&e��`g&Kى�x���x�yG"����>/��}�h=��ۅ6�^�e!�����a4C���q7���E�9;��P�?K5����bW�#��˰-�.���09Ec���)~L� ?B�U�L�d�+�Z*�U�$&\�5�D�q�?Y��2��݇+ ��To�q�2� 8K����Љ��N�{����	���84#��<��G�x�bZ�<Gv7"(ڲF!��8���ӈ:l=kڶث�Qw`���s�@��K�&P��Ʃ���4��qI�kۘIw�=�;a��,_�L�LYP��$#f�����E]��_�C�⯍9|���@��ݮ��NA�zj�<���o>�.�� ����>; ��闼[���t�f�ާp�ޝ-G���f�,OT��Yܦ�~>�>�ME�|����a⏁�h:s�:%�F��R��Q� TI�tmn�%��a��CAc`#E��3��qģ�+`C92j*rY�c7��Fu�|�D���T�-�Av��˓���A�YH�i��8�B"#ઉ�S,��$�!�':�Bȓ��{��������N�.��6����M�Bs�$�Zl�� ;��.���7�Z��_�������"���x(~x�u�3!R��I��M�T�;��i�,���PvT੗���c��q�nW(H-�����^s+y�~����J�^X�p�{�~H��虸�S�ދ���,���򧽙�F����.����V��?fDҘ#���g� �A�-�p��~�(�����]i�Q�9��!@��Beҏ��"�iSa��R�̀V�0�3��^�in
��k[7,1��J�n2M��r�S�N���)gI�� ���m(;Q��f�e��u9�Ȟ.,�t�/ӛ[�lI��Bim�N�s.�MĚ�����p�۩��V悞�����Rr�ww�J�E�;?�tZFk�V��R�XG1 ؛�]�B5� Ի��� h.Ҥ���	��
���}�մ�8��|����W��'���ʀ����%;�άl�Z<(���l����i�S�����h}��P��38�F��jW?DƔ�QQ^�+��a�a��9��El;���A��r�G��Ľiڲ[3Ƞ����"Wxq�����J@ 9���`	i4p����s{2T�/7���uE�v��=�;F���!<�ŝ6���K��~X�m�wx���~���( L9���χ6N-rj��e2�c�ұ$���e���[k�f7��
=O�Be[&�k��rХ��ˠ��?(Dn��uQkA�n*����_1��98Ɲ8g���v����*�8�t�\�Ha`7��Y#W���`��/y�]9�ޘ�����#��#�UTY��W�T���Jo���(ɗX���84��_I���xcH� �%�S0��-��B{O��a�����h,Ig������������
�/�I���K�H꒙vb_���`�]V�����k�u눏������y��*������m��-�qB��-��L.�J��Q����ʶ�*Bi��T;ԯ�zs���LOu�gJ��[�>�&k��5�i�4���jIx�/�X�'(�M�{"� �9B���?� �9U�%؀�:��/�&u��~⦵�hU����o8q���|mS�����o���c�[{|�z?*�j�0 㢥�}�y_9��u��z�:˧wK�-�f�.�n��f^�4m�Z�[�7pc\P����3I�Ll�?�=��� �{�h/��G!�,���?[;��3�K�kI�'❐���)g�"���ބ6���c�Z��s�=��Wq��p��=�������0:y��1�Jr"�6�A561�h+�ZRV�>힩�'|� c�OT��R�9���4$Y�ĪoT����͉,eZ���ǔ�y��h�B��5�Q���:���u5_�8���7�OSNR4��܆�z��� �#�X�K*���]n���6��>Js��tҜ�'�C�O֞4)����?)�ذA���\���ޓ�J��$������4�?�II3�������3�$��~J�c��4��e��=IQ����vIU�"~�[Y1)DOy�
��H�zI/�bCZ0������4�㙝��#��b�s�����[_W4,�+��U@�M���m��P�2��pq�AV;�V�� iT��8�O5�4J>
5�[���)w�������U/�h�S���Q���$�TF� U4�`{J������߃��%& ���843,�YXX��Ti�*��O(v4�t�d��P��@cPk�K���N����W��r.t7�4r�ƒ	mV�Ò��ŕ��ͦ�.���C��$�5�y��@�}l�J��I��{x�	"5���0���,�?	��f�y�^��o�S�A���X[5j����F�����-s_ ��s�g��z#��E���9�G����
n��ɕ��{?a<Ӥ�������4Yy���sÛ(Һ��D�@����Y݁_���&�vNJ$
ě�u��M�R���Qa��\�T�H���9?�|��W��vH�L)�"�Щ� -WzD�ZL0p��0u��N�LZ�!���"��=3�i��e�dnJ���������}_ϵ>��we�{�
?��B}���y�8�&�l�O`gL9��3i��?,��s�@�v��
s��t8�x�M��?
��r�����H! ��b��3y0?�H�O�&G��p�\)?#�$靈ە�S\�N�O{/�׽n�P־`�,�5ty�����2�Í�l�8H�0*M'�b�'Ϟ���r:ݒ��Mg0��$
!)�5K�Tt&.(-<�U����\;U@)oF�o���f�Hr�5$wG0���ɏI�ד
����|
�<]ނ
��-cy?o�/SH�6�0p��
G����ߪ{��$,@í�����K^�O��pE���3��͕
���F7�R�����V�HO��-�_�%����t߅��|�;�����Z9Dw�r����������h�IV��(��\���1~��7���ElP۞�"�o��I�ޒ/r��3�q���X��c<��7o�]�kfU����|S%�X׻[��M�C�����V��d���i�k0���uƟ��0Z�l����=3��xF�Bl�\ܒy��S'�R����T�&n1��8�����9\]����棨�xRsf5۾�4#݄'������?�/�@{�+��Tu�ͰO���u��ׄ�fI��*�~�]���T7/�T���rvG�n;�mBx�򇏬�g1�Kx���r�?bX�|�}E���&F`M��@���Y��>��#PP�z���1koK5H�a��~�\��P�F@��
�y�@^��r��E3O)w׷%�_�����fc�ʰ�
�~$Xhaa�3{I�P9�ټܮ�S��q�@���ku�2ƽ�f_4�T�m��s2�$q�K�ݿ�;Ll��V�D&J���Qʩ�q&x��(b�a�|��~�J���J�'���/��|%��6�!��U�r�7 s�~��@�:j��ڐ�"B��y�Oo^$��f��!�yM؝��>�,���jv٭'��P��c0�)���n 3�tFwy�,�:�>��:X���k�U�,�@J�N~��_���Q �A��	q�Zz��|�f�*_��Y�2x8n�����E����O�˾�����Ns�V��e��8,�>��}3���%��gAǟ���e��vܟ���Q,��#��ܷp��ky�LQ�E&~o+��8Lb�Mw�sǞ���݁�4Q�
E�����3�ї#��.է@X�����F{B��jo�#0�FbP�b��~��Xp��Y"�ey�
\�@vRF�L�:�k�<�<HT(���Ԧ 6Ő���:攠֦L������ANc����/� ����[�y�	ӛ,���X��0w"Y�]��R�/�.]��i����o����l^ק�>�'h������5�p����@�R��«���?�1�~�M�t�X\�[�}��%��v��y�I�&�f��E�:�=���_��u�;���v��Z����l�=o�#i[�E|��8ޝ��`	��r�L4�쌃)\EЮ����Yp�R�S��4h�<��o�1����#�u�̺o��9Xꬋ0Шq23٠e�)�I���E	�3Z����vְ
"ɜp!��EO�<A>Fm�F�7}�%�!<��-��b�͑��/~�u6�W[t��3��.8�6��&5�d��Ѿ}h{|����v�$���d��Y�����}#���l6-�ZT/�G�1�5p�.�ès&��X�!���2	���POmZ��|�d��}�]𬖏��;�l\j:R����8���3�V�
�\t+�1�y�_;�¬cC��a��Ͽ��/��f 9�b)����G<�u�������%2��px\�۠�n�'a��1 26�PU3&%�������s5�We3�	\ȆAԗ[A}?�߄n�2V���Z�p4�>k�K��M��\E�}yE��������{�F{�Y��'���&Ze�Q2;G�0+����JiPe5tA�Dt��X|W�;/o6��5���ź�U$z[R{���8I�T��~>Ϛ�QR��~I�T),)TOQ�$�Wa��im��>����	�_󋿁H�����}�ȫCj/ܴ.U5�EPޤ_�SLaڤ���_ţ����>��_j��B�X!�xb�����P��m���`b��h��6��X2)���>n���e�����)G茤�� �*���7���m1�� �uv���Y�j���>����>��I��t����T��c��:J�5�I14��i��I�W�J#~(ǩف�B�cu��Hd Guc�t�z����)$���z��\�6��]���4��mt ?>�y�꿽z�C�@.�7ʄzT���m��	+ة ���ň�o�6��Q�ev�ρ�����顈��n�卨	�v����d7HI��4OB�1!��^hV��Bt��c�٣g��f�X6�-/Y��w��_ٛNea�-��8Ù��q\a�9����ʖX�y��ԙhLY��y6�;��|�c�-���*���+Wm��|R{J�d�/����˔�ύ$�~�<?�ㄤk����h8n$�8�����D%
����a�vc9��,�~��w ����I�D\�����R=* ӌC���?N��x�K�\����2��� ���`�,�}Ƹ�ȣ��L��f
o�L��0���X�Q�C��7��{�L���cf}��(C>[���_u�2���T ����Q�9�ZO	8�JaG�k���9�42f�-�Q�� �P���I�JѪ�b���R�z�oTI��$N*�|TZ9���c��Rp��Eh*���?{.��8��(P��S��6V�7�|�^��S�hC�e��),�
6������JC
�l���UB�H�;B�.$2'm�50��=�K#_ǹ��l�{Ӧ� �����΋��{�R�tU�xI1 W�d�X��PW�f�n[r�q-���LFU���i�!��T����86B�5�ȩ"������B�Φ� 9�[�u4vT{
��x��9�<�%��������sz�C�H�p���q?����.O4���4<��
��*[<�(�f?�9�������ҧ
/�p�v�f��s��FJWS���gt~�{ڭ�zK���~��|�da�	��-�j��r�ܖ�o��[�ɬ%U;��V;\W��x���@~�~G�?����V��a��<i�3Z��A�r�s)��9T�C�oy%�#<�<��JHJݰ��x����>���8�
����T\�Q7���c��B�.�Ka�?�W�$�����F���:���g5�j�Ϙ1�<�#-hu�q<�Z>
����9����������[fUK�6U���<�����.�_.i�9FW��4������S�p��O�(���(2@��`T�ܳ!�k��4�7�"�ͽ�2�,���E������[��Q����Ȥl���:�Y�|F����Z<sr���USe�Y�Sq��9Rb�E��YL��ݪg�6I�vj�ҾxDp������g���X�e
P�k (�ДQ���I?�yڐ1W�4w?TY惔�I��rS����	�M�"k5� ���r��R��5Q$��09�?�hd�b֪��v-��bҦ��,)|ZqL�p�)�'U�ڦ3����E�x�����=h������n���7'[���:[�d��a����0�~��p���1�s����+�����E,�9a��f�z-z�^|:˟'"��k�f�"d1�ci��~�,�OH�~�t!	�`a�b0�Pߘj���: ,r_c$��� 4�ǵp�<��tX�1W-���w�Q��S` cvtA�=���b���^��9�`\����L�MU�pw@ry���rS5i�+^אա���>@�|�ߧ��Fb��2�qξSow�Jsʷ�v�����6��qMJ�mN��
�4ܼk�]��6�T_0�GP.�@/��gJ�*=l��|f>�
d��+lcu�S�"�;��Z�S��A��
ˍ�ΰ�R�Ru� JҡƩޭQÕ��4��@>i�����fi]Z����L��R�}yb�]��OVx��0el7_���~�RV�}�)���LFFH��*"P"{�#�xQv���j�3�����O���{_�=�C>Vo|"�6� ��ET�1Zls6�Q�{ᣀ�J�u���w! �m�����B�s�D���7V�����w�,�\�}�Uv��p�Vn�q�>��G�
�����[��:�������d�ӯg͌����2����ܔ�}Tl����h3Q�@�q�""Z�e엀z��1���^��v�������9W�/�)O#h�SJ�V=*P]���G(�B�{��-՟Hh�0l��hO"p��� �C�f�Θ��P�b�pƯ�T�P��4���0_̓�z�$q8z�ӄOB"�A����9N�lA������5h <��!���m�gJI�*0*�O���#�������s
���&����=S�-� !���i�7=,��"�EP���9th��4������s�Ei1j�sX����~����b�q\AX"�Z"�D����dM���������������F؂�y�bZC^�e,�?q�@�|��Ml?�5���r�{��#i�[��^+���|�G�{��K�}��.!�=�[��*�m����
�a�
��"�7�M�Big���9���1]E�{�͗�N7�L;+_Ht����|�H��:c�j��G��L�Ju������a�@��(A��P[�4X����9 !�e�08�K�>�d<r٤:�e�	��;bwD����aU�����BVG��4p��i�z����nUςJ�bQJ���qG�����?-��*���9�h��h\��p�ؗ��?r�o��3�y�#y�QZ?}PX
xD�Fط��e������"gxHk����b��ݻ�X��j����1�ˆmَU��~�RD��E�[r�b�L2�XF��"�KOmm��m��6/�5o��g����E���Rd�����w �B����{Z���mx�k��JT�8��s(c��'�F�O�|�����6x��b�x7svP?!%��(D���$㡡/��ڋ��U��ێ��D�G��������c1aX,�:��L����\@x |�Zqj�d ���T�v��{�i[~-9�D����r3�MM�4����ܦm�O,"���ne�a5!5��8T�@��3����i}|��Nʶ��ɋ��ܙ�O!�)��d�̗f������^2Օ�j����V�8�5פ��%�s��\ %�	er<a�Dm�6�OCz�3��Þ-��s�����Ȝ�\)�_���v���X���o%��	�N�Ꮌ���C A�����.w1�
E�?j+��	��)�Y ��t �ݙ,s�6�"~�ƽs21�j R����-_=ZG�b���s�s��
���x�%�P�/���,��ֿG��g��u(��B�W�v$F��f�F#�1r&�����%�/u��ۢ���I�$x��>6��<05K�j��Bɻ���
|���͆�,1߳��
�c[2Q|�ДN����j�1&���>�Ӑ�0@���?9�p��ӫ��4����w��y���L-ծr��
��h�(�H�"'�S�����5�U��\�{<��w��1>�Ӌ4{I��r�t�d;z��]��������KT�L�����n!��LC)Xqh27�hXçQӷF�?�-]#|�ʉMVf��0ޡWѤ5�N��ط�� g`��\���/%5]�F��Q�+����@Y�+�tF�.w�,`���z�3áe�X#	��^|��	�;~^va��"Re��9xmʕ=��lw\ձ«k�0�e����f�L��ݭ�&��-��@�J��w`��5X���Z�O!�-OP |,����������6n9��fy��<�~%Z5@�l�KN]��Cr��%�F��h�+��U��@e�B�ķ�ѫ3��Ax����\憩.��+��M��?!��4��VG�;�ȇGv#��{�3j�:�l^F1d_��mB̒]�|���v�&H���O?�b�b-�>�A^�9�d��Ѽ������@C�l����$�*5�+�ݟxW��"�Ӛz��P�ŔS�1n�*�΃l�-���g%�o��w"�N>���9|�|4a�0Ł�_o��t�l�٢���N�b$ĺ�_��h��؃kcT+y��0O��w��3-��I"AzTfҎ�8��^�IP��lT-�*��_lK[�n���&��R�ߣ��V() ��%ě����S=�������8����/-���
��>Ĝ�R2g2YE��ak8ʝ�@ Ù ��������$l!T��I��M�衪fLm�Z"�R�l���|���0wy��[C��WIm2��9�2�;�{��4�U�I���Xq�Q�vNL�G����np�kŴ��"/Ԕ˗�᜔`\�BI\N�g�Î�v2��w޼ի&�n��O���Y(�� #�7���J��m�b�T��Ҙ"5��i��!M�
>���@F{�Y�m�=��&Y�}�Jv#~!�����[�頺�U�>�ni ����8�;�#)��<�i
5DXJ���h�cx��AoZZjdk�D+t$�YG"��@��c�s�?�	���<5�� 6 =3잓x(ˡ5��WN����`4ͩ7c�(�໲��؎��Ne�%-S������� p�G��tWf���,���+R�MSo8ɮ4��� ��Ԩɮ9�8n��Rܠ�l˕u�:�^�-{@�e<�8���N�Ӝ�<�0���^|���p�<M�%^�E۹��Q|��+����P�-E�4�����c`��CS�+|��j�Y7�>�֡ŜAT*�O���w����I�3�p���"f����0c�N�7n����5�z�\��T����:���x�s�h:�vn,��KA�P��5
MB�a�a}����#�\�=�s����mj[^����6h��o�#�B[�>�J�����ةS詗�j0��7`HW�BNG��L� ���q���s�(�R	�lE��^���0���s|h���wf�'4[�S�K0;g������cm��wnɋ�|��t\{��h%�=mP_��
~4)�r+�)Ҥ�M0Է�+m����#��C�p�@�G��!�����<(2��g��E�(����]����C�Y�b(��$:f�o�
��؆Dgh�h�L��ܔ���U���mp��^�>5�'��#���j,����T�c�c��d�A��s3�SLg�9��Y㮓,'���d��ꢩO�O���}��mۏ\��{;���ncj�W�:FBs&���ȵ>d��1(]�i��;u�O1�� \������$�'�4���cv��k7@w�̇���S�\ɘ��?-��r~�󛅣�Gf�8G���6~U�q�v��F�Sn#�Eɺr��*��F�vz�T9�=�rs��D`�G�R���nڶ�>:)�vؠ�$,a���q��?��M!^iH�(�K���7s���P�s��2���P�G���Q�׺�	YC��M�n`�ÛѨ�(��[?����%��W&�ӏ�$�$���(Ѹ��ˑ���m9v:\2����`Qo������(��*U-�jj�W�]ᄠTj��t����g\I^<![D�/��IN @�(��?�AP&�^�1�|%Hߺ*�%���9����T^�J_fo����+��-�����ą����g��;u�����!��|iym�n�������1�;�jDc7GS�HdU���s��5-#�+�1db��!��"~�O������m=��i�5G\rZh8�qe�;�-�Rj�gfJ���f�5)0;�]".�"��Y6r���ʁ;`J�:���5��춴J�L�x�w׼�sk���y�`�z�ҒD����^�����I�(�M"C��Q��,9�����{9>t���.1����h��EK!	����?I6q�ʸlb�O*�NcNr�'pE.�'x���#G�ӡ3-�Y@�D�F/3C�|�hQ�[�E�1��v,P��O�j�ΨfҚ߅|�F�&����/�)�)�a�m{�Re/aB+�&c��k!�R>B��R�?��p՟n{�[�iq�_���W��`-7���R���Xb� �EA������!3MB��c����O�@��g���0bTA�M�mF�6��9���n~]\x����[�#4�����);W��:��������Oiߛ��x+Y��wM1���D�ph������^w*�Cg��2짰~�K��:@�?��^_E�����
p�� T�-ٝ�<�Z�r�����\�r�~ ds��Q/�K�0�FZX��]�9��\�r
	$z���Li�ۧbL'��j��6&��@.���� 7�<�4�A\NĲ�gⳅ���]�R�'+Fy�ʡ Άj@��M�¹��H1����Θڊ�%��~����|"H��Ar�!��Ӂ� ��ϡ
���-3q)���IѺ1'��n��t�+7����X]C1��Ŵj��2C�����ƅN]Ys� ��#��ի.knt[�l��
�\d��-��ˤ�xދ����iPmT�܂���|$l98f�o�������O���juǈ �1:V��ܡ�+'ys�t����#�C9��_�Z�d<>�@����PE�j7pV��X���f��F�G�h�5�~D�6�n�����G�5�P<� ������-��S��,xk��X�zP�c���뽘��w�A��ݝ��T5�8���o��SV�Ǿ^]��eU�W,�LS�5����u}����8��F�'rg5T�{��]�鑉������Z�`Al~��of����L�9�����p �K�В
�5�zA� ~�$��]���v,Oy$U�'|�>�9�C�`eg$��X�M/|q��6�K�}l��}<�}���W@�&���A��QR�
�{>��b/#~�7E�',u��cYo�r�����pR�
.9�L��r��KN�*\b��sz�5��>������� �k�������>��	�N�ژo�@�+Q�,g�����.�`���������s�� �����m��z\Ё'/So�K_	K�4/�e�,G��6�����wMk���}�������a'�:#�+�)u���!s�&�X�cɫ�i6�b��xS�1B&͇#UFt�&�D�;��j��p�c�tgbV�SOnv0�[�W)��/���k� b����y�Ǐrf ��j ~��~:i��R9Nxc�N_�4G�Z�s�+-����N�`�5�:�����d����P�f,�B���'������`u����^�)w�� ��������q��כ�4�wq���9v�#���]���ʢe�x�ǀ���f�� W��j�>\��|�*�+�"�!�XT�����ໆ���*oK��=��b��h�����V�ɪ���������&}�р�bt�4��If_����1}�o&�V��f������v6�TX�5�B�^r]���ZJ���&q�)�y�:����K�}�N$~V��ǳH����ׇ(�j<8.��O���Ro��za�t9����5f�q��*�����|oǆi-Ĕк��Ѷ~<@�O�VBdT��0^�ŇdZ w�bJf���6UG�Z@l�./֞��� ×��
��^�Q8,��y.B$c8ǳ�[R� ���y��Lk?��;����Ƚj� �;��H��:��J	�{V.�����mD�4i�.�j�27�lJ��+�;y�I��oh�校ɀP��ͮ3�Uñ'c:�[���pz�F�l�BBw�e�<�q�t˧dd8$�
�c�G��_����%�~o���R����U�멪s�O�o�P�4Q��<��y�y�Zm\�y T�Q�=�X�MP0�D�6���>O0#�9L�s���16�����>�� �@F5"1�ګ
��ڒ�b	*�H�GV�s"�,����b����H��J;<�코�q8�
r�ǧh3�|�O)n������k8$��ʼ����shK�݊+' ;�o�:��t�#1�����G�#��g���2��߷ �?>�t�%�Bp���I_�xI�YO*#oT._�Ü�-3u���Q#h:�A�� T� qǟ�(� 2���5ޖN�KO�A�n��=����P�v�'��|S�BL�z63�f��Vz
jD(�$1�����˟�<{��q	�R�W��o��j��[9/�at��[P�]�h��ҏ�u�>�c�H��H�f��<?��Ø'hM��DTn)8�4�7ឿ��;2�Q��
}�mT]��i/ZL}�ص��os6��%<iȁ�N�s��׆��7�^"�d��
��%m�V�QC���Z��g��l�I�X�f^EbA�[MԶ�B��b��G8;]��r��oYr�;z�KAMYH�@�H��á�uݞ�i�#Q�4����Z@����=Ԝ�ŧ��o-����V���<{-G��W���
���8.a�;����E�Wv�!��jd^jK�<��BN�$"k�2��G?4�}M��϶و(�	��a�/���7Y�<<�V�q�(6V�5߯r�C$�=�*�H�\�ӹ)唳y4BR�.�TeM��8��������8��,Nw��u6&�. 5���2f�D6\uH����2����75�� N�[z��3���lsA��L�SR��}/ �h2��g�D&Y�A�kț�q<n���P2&:�.!U>���Vs�����Wv�n�+��w���Ӌ�M��1S-V=8>��BG���:Q�ѫ����{A��O��=�A��/'�$��>����U[fnN��G�B�`��Q�4w��3%�'�D�J;n\\���tvm������Y�(�l�%�&�e#Y%���Ht��l���Mc x�h��Y����r�U}��^�d�B���Ӏ����7e�x}�ƥl�(���⠧b�~�#�h1���M<��U0J���JgB�hXJ�/ �wѸz�xZ�w;.� RՃ��u7�yd��e>�����O��=�Q�'k��Y4۬*ѵ�u�2t�g���
� b��2��M"^^V�����kR �y�I$
�a�3����Y��$�V�w��W�1.M"�!l�W��w�Q����u.��]G���GC�3&��b�I�"�<<j$E����m�;:�M��T���zo�m ��Rʢ5�hӉ�fv�7up���C�~KS��M�j�U����^����2���kQlyIЎ��7���0�~��z�a^�'E��Q��L�w/k����P�)�i��8�'�]XS ���jStK����4B�
TM�dR� ��� �_�)1�*<n��v�m���J�3��!�j�Gr<8H���9۾����~��` �<�����dI�<�T�>�|B���TGsgss[�A�u�o.��:�uȸLX	F�{�ԡ�dw~�z����O�5�ѱN�W�����s?�Wm����mn]`�S�T���K
�D���E�zn�kI�y��4������Q��1����g���}>;�)ԍ����R��a��(?}=�Q5�8J�+��$G���iΙ7�+h,f(��(����P6������
5�Zk4v�Z���,S!p����"W��`��h*a6C�L)���)Lh{���J��ucKQ<|�R�#l�{q�DeJm*D���O�}��-�� _*2ǚ0EO���֊�3�5�D*j�|`?ں��	?�����t�8��Zh�1
��X�Ռ\���l=���ȞK
{O}CN,~��*�Ü�ē��'�l��|�q���=�7;��> �����+|Ǥ�T�ƚ<��@�04IX�c\��I��"�C:�3���L�FXEê�c�뛃w긽��y�l�r毢���j�&h��#�";�G��AI*�"�F�粖�h?��gr�Hw8������L�h�>�է �GA�XE�����媌�2�r+��*���?�����m���� ���4��	��
r���gܔWX�A���,A��w,�WG<s��Ch�`1��Y�F��>]=P��L�M�uAndpiz��5[�E!�H�e�(Q�c�~���Kuo��1B������՚�a�Z�m�6��{h$�z����!�uo�⿉$�P�gI��b�=����ea�vzW�
j��i(�*����+�c�ͱ���zSGFY�7�k�:kϹ���o���;z�;2��:��ȁ��|����(����3	���YZ얾rt�$_�� JoV�G꣐�����]\y�V�q��&u�=��N�.h&��\�Ļ���~a0"�av.t��@����	����=�PN3�j$'��4�%��c���aA2f�)� ���L5����Q̼=���A��H*z�Q�r>չT��m���Av-������w4ñ�&n�\j���c6D k����~p������k��?�>J0�oYLSW^��ыm=�b^�:��`R%�q
�!��}*D����|��bTPz�rV�<��㇡]�[USw�"ᔄ���z\����y'K��M��-(SF��6ϴRyNe&Ѽ4"y�.3z\�����+k�П�7��4#SFx��ť+�u�yNNgU��K<�S���q{v��F\v��[r����4�0����v��Ba��*�l�z��k2���È�_>V�g�W����#�ER���?E��9�կ�g^�V��H:�d>U�׬�4�ڇ#�����MdV�+�{� xI�8P�N2��ʠd��A}nJ��5�ƴ���Q�+��׌WV8�^6�6(x�oOL�o��	G�S�>�"��r�"�d,��[�	�~�}��?P܏�۟)�E����Hs(��胊���ͩpg?+�%l�F��������w�,_�%z:�ҞVb@�D極].�|2ѿp/ۛb mNΫ�=�l$*�g�|���l����}q�J���V� &�=zl�,qoi�z�?i}�ũ"7����َg1��Sf����}@�-4���>����*��:�t�[2r�Zi�)�
|�+��/�&tQi��B ��c�Vq@Kɪp��T_�zw괄e�&�z<��=?�mk�DD�����s��ϵ�B�&��g��]+1W�ò�̌ݏ�s���K��2����|��*�v;������8�j�������k$��yv��G��奎�:�E�m�+�����Mm+"<���(�6��U!i7��=�z��X+�O� "�@Ҥ�Q}��y��q�����W̘�ʽ&��g�pw�>�t�r3jU������4L�{���UY�^xh�����Z��W�S��XTR�-мZN��D]����k�.�N��JN�hf*��� Iq�����H�fq�w_k vwIx������+�=�˪\�(��"�M��DW��W2t<�C�1�(�k��J����}K�J�ήL���'��>A��D麙�A���̪t��v*� wjc�u�]0�]ZT��gt����C�5å�	�/��q����#��;������m3
�+�~�����ҵ�78cĻT��mX���f�;�E�փ� �N�2�9��ܦ�T��ܵ@���3�q; ��>澞�\��������'px�Ut}]��5٦pe(� T�5�6���+IS�z D�" �XiNE�	��q�T�~��%���"@l\�ΜAc(��6�*gR��bH�O�C��z�d��捣όs���=�1�r�I��~�6HO��&��H�f��R�p>��].yu��3���`������u�,����k�X�*b,�/�Q���ߒ͕l���`cJ�mV\5|uN��z�i������:��-�F)V��7]'�u��.q�[ܾB:����>$�fN�� �%l�Q+�x�II��T*YbS#�����S�o�]���K �ܩޑSo�D4�jdD���-Љ��r<��&4�;��w���ژ ��8�,m�o�_��lQ�����8�D% �5���2 5�̬��B�$[�pztdT;d��(L��.w�5�h��.#��u��u�l%l(l��D��)��}��Y�i��_(�Wg��$���~�	(�/���UYM;��� ���iI��vSD��� ֤�0�$1�̏v^�����8��^�I ���d+ݰ�+����ۥ5ζS)�]�f\���JBYf9��w V}X�V�b�����wB�� 
��o&�Y߆$��v�
1���6�ϋ��I�2�ۼ��|�Xbb�n��I��<��	�ͨ<q��5[>R�K�ԇp�1��>������q�W���r ��`  $�����s)�wj�\�Q���"��s��y ��(���d����E�����ח�O>	�:��.eC�=�xqb�4�H�9' ��P���wEq�>?�[)��
��b2g 0ό^]ES�ucDdrv����,Hy��[������3͍R���Mӑw�{�H�ߑ9�rF�F�x��'<��&����&��Yf7Σk<1V��
�(��*2l��	#�ԙ�Z�vI�-G�����v^�$m�D�-9�H���,�#�Ok�4����Д���*�=�v��DՖ@�b���*|5���B�!��&73�^F��z*��_�!��Q���?��9W�Y=���s]�!��Έ���Ada.�}���t�,�Ԁ��M�N{�d�.���;b�U�{A�ܸ��

Ǧ���eo�B��Z�2M)�7�(q��O� -���ykX�#}�dc�J���5��i�1 ��h�I/���{�v�u��@x��-�K-ٸ����e��e'�G�����ZK�,K?F�l��l�l>ٙ��ͥ������X
Q�Z��e"��,K�(���_�k4��J�z\������(����� �ղ$4c�p���A��;p���{�|��ݤp�j��T��ERx�&��=�Ι���U�Y��Z�Ga��~�WEOF^�El��(�}��=@����"���?�"]�'8����̖�{�^������}B�GwXJGWv�*i'��}��&Le�'3�������<!,���Բ�ˊ4�=!���N�x�mv�Ú���yu��q�*��꿨n\�/E��W��lT���Л�vy�aJ�����Nn���!t�Y��,M+�]��3�!Ȏ��������{�lE�T*|��H	L������GS-ޞ&���{1�P�A&�V�=��M�A�>R\�� �cm~\ZU��L��a�s�wf��:�Ϣ@h0-<H�r%���y1��K�O  �T�7�Mx)��=��y\�Xjx�Å&�7Q��C�ݰ�V���P��\�-�1�o/Q�?� �ח��V�����b��߽�&�3����z�Lve�p\��/5����aW��w��g��I��]�=��u������yx�<�+mF�c�����4N�~�bx�|��?'3AT�D�^_M쑃IT:�Gy<�"�h6�̀@�	�/���\�?(,�1$lG�6<c�V!�hbB���b�.�6���2����_��mU>����t=m�E�����̸��	���J����va���An��Q�����q����T-���$z̏^�:v+@��p�
׮ת�8�ޗ"��om���s� ����軘ዂ���H�,�h��֡"��,���-�b-�7�,�c�V�z�@���/�)Ej�O�+����<��҉�1�=L�<����Tb��["ۻ��T���Px-o)��Rz|�8@!�U�#�r��A��ӟ=$xQ��B}	%�D���	�Q������4S��$����t;�~����v�ɴ�Ӭ�B���*��P%Px�ӻ���L�t�ޗs��@#�&��k�pd�]����(8�s�z��"��`$�p�y!Je�v�~�L����g2��0��>,���Q���͡Udu�4������L�+i�t����f��(�B������� ���C�.H�>�i�9�?����m=Q#a$Z�+�b":�����y{Jg���A��K���~�Q/3.�O�%�J��l�����	h+7�N�Jq�"�qQN�s=�A�؂�ok~�G�	���/����ؚH�/��x�j�ש<ѵ>߶���pi�Z�D�s>h!�X6<s6�ؤ9�VY�&�(S�����'�N��@���
Nr0Ɏ���T:<�R^BV
��b�F,�3fvݷM7��b*�%�k{��!>~�a�\���X4�̭r����5j�5ݱ��Q'�)@���En�\��"�ɤ��;��q���i�z��fr�OQ����������M:TB���H%M[���ݣs�ɖ�&j��K�1&�|2��wd��j:�ݪ��o���,�4��bg[Bc���[���"޸�;��'��]+���*��+��8����F�`N�|8�$,��BbA�3sd|�*��ĝ���]�-��{ה����	�9�lp[�0!��q�x珯׾d'��(���6-�A�FR�JTk��uj#;^��^�~��� �"\�R���xKC�_;��|����,���1Rb�$���B�)��	$�K����r�/���^���f��T&Yb�6�.��͹0���Sg`Q����X�{�*Ϻ�/@*o�h�I�4!�e�lI����!�u.����'zk7��f�=��-&q�Hw��f�>��R�)ѧ�~�����]uR�B���	τ�2�p���6W�,N8��MT��h�����i1�<�.$K���t�o�1·Hp���a�Y��|ŧ�m���*��!��'�v{���fB�������4~��p,��������Y�]��8*iqK���zȷe~����+� ���a�1'���,�\t^+�5j>��&b?Y'�#`h2�$�
�oXH�Tݮ�۲J�9��1�WM�,Q��<m�8��ֻ����7� ���l/7ѩI�џ�B�>�)䙤l�\c��������uO��:L,���~��>	��C��/B�>v��W)���?�uA�C�$����OJ��#s|�^z~�\T��.�u���"��d���_��s>"�vקۚ��|�3�hT�]4�l*u@�ݪ�)3ѷ�S/�P(Lc4P�!����50���2���A����/��>g�T����B'9�q�_���� h{	E��������F��9z�,*�2Y}�O̩�m��5�ۺwgHQ2)����+7&��y��5��Y���$�a+w�)D��0����{m�!#ԗc�����a��Y���-���mT�Ȓ�A(��沫���&��4lgD?|K�P%;u�HNs;�W��3�i��/�U�7�ݵ�oL���2�ͭ��Ҵ�L�h,.�%�?.�'�BH�0� �h�^V�<���q��+@ �_Z����[�Z��й��LO�f��A�(��e'��P�9�7��f���0�p�L_��FP_����*�c��x��°Ʋ�v���9��X���^�l��Z�1|f�xCzz0\����[��D��BD���Xk���F�N����9��|��I��ms��U���&[IIp�mql�.h��eP��o=�8�,}ݛ<����u�0C)�r������M����f��ۆ6�VB��������Y6�B]|���I?�~dZ��=4���</N���s�>F�<&��a�{E$����as�X7�O�L���e|N���8��N�Å��bk��[�+� �=�FNS��dHe����{��(�wH\�rb-Gp���Y��XsK�l`�ٸ��N=�� �7b*U�+_$�0>��1h=��9�j��������L+�y��i]+H�l��fŃ5Y+#��Ŧ�`;A�	+�3���J.�fц5���g��2.��Τ��0y��K)��"������տ�۽ohf'J)�XWZ.��.5��pa-u��hm�.ҕݴx1�~�Ig�![7@_� kwhm��)����JG*�&k�4T�Iɴ.�K����qo�m�S��&��p{���Dià�#�`��v���f������=�Mp���ϒW�}��1�`�B��I���iwZ�z���7�9�����)�j�7`(�SiD.i7��r$�a$̯�	�|/y�����D�|/�b߿5��I7��g��U|[6����Ls�[���fJ���0��iE�u���UI$�_�U�U��8�X���9~���[ZT^K9�G���~V�H�w���|_s��n���uQ9���t�VF|��ժ؅N��t�\�lL4m���4b���(J�ߺ�'��w��ړ��?Vr���XӺ�a�봒���8�"y4�}����3��+��F���E��E$�T�$�M瑅"���9A͉v��0��[#
X�'�5�9<���Z^*�Rh��
���EN�!������}�����V�zM aNY���l��N�/6�)t;��B.����Z�H���bv8�C=�ޮ!Ƣ�O}�2�����>,���xb��<�x��`_	��7*񍞀�#?�ժ�N�9Z&�K�bR��M]�k��%]p�D���˴ٰn#K�d�2޼8��ͩU'9ʸ���Zq,کy��~[h�G�-;u����\H
n�P����ԪwJ�z�n4�������������$���Y����ܙEll CHoV O�'h�A� �6�4�lJ%szfx�[G��S%.a��8��h��2�H���=Y=�(z�q�����b�o���d�:��d�5�6�ėg�C�Zw+��'����Pw����,�nsd�L4���YөY�@��۩�;Gxt-��Y�@�Ck�����md>�,���� �cDfu���xd�p�H~4п�
@q�}=0tK|��X�D���nc��f=k!u��-w��L2j�y��&?F]������;m!�A����\�p�6MK��d Q�u��	JBgX����&�T%��:��!GhWI���2���8r�=�CE�0��v�(��t���Y,cm���~2sq�qZ[sADXSݨ%�T
ok�1'!3Yެ����v��}ˣ�eM�s/N�����X'���D>�b�Ov�	���dz���,��|7�ܠ�}�v�~����5�F��ʬ��/�B��	@��{���w	�(w@\��E�es�A�<Y���3#dF�x�H:��s�n�<����:��}r��:��π�ݸ��Ԙ�uʾ��k$G�{�z�I45��4V��_~އHA͙�nj��1��֬��CvW���m�������av��ō>�����4�5�}}��`{���0PGb�S�ٲ趨o=O��>�V�o��ig�S�	�$1&CF����::�ڇJ�RW@ҙf�\ow��F�|���]q���4�R���@6��)�A�dw�C��+���K�3@���NEs�}r{����_��p�+��H�e�O�m_�j�egu��L��5e�Ro
˴�W����Ar�J�d)樚�`@�T�e)�I�%�Y����iw���D��qұo_B�H����r��F�9mj�]��p3�,$�{����0���Y<L��!a�yY����3�P���/Yt��D��6>�9�=|<�i���P�Y샄����LM�<�Yh�Z7� "�S���F��.<f�Ys����57%�f��9~����h�>4S�l
�%��*�xLYfP	湉=a����d�U�v�oPS����	�<��{�s?\����\���U�_�i:�w��;$�h#����M��j�p!��v�lJ�t�m+jo�+"�Mҫ�P�}��ϻ'�&1�iȡ����9��&ۄ<��^���l���	�̆|�	�t���F��V?��(:��Y�1����-�=�C�//�]��z=��1��H��a�i{}ђ_{y�@��Y�Ձ{�N�U�N���,'��hL�fm�:m�N*v��VJ�@K��<ut��b�/��4��P��(��A@'{tM1��y�:�1=�pR�%��^��b���m�|�u�d���[���B�ubBm���
sA��ͅF6YI�`G*�cq�7���ե���4�-�	Zr�P���.�h/��,�T�gbK�N�P8�'��X&n0dn5vР:��@&WP������[W���/��������� ��V��л<w3��Ά�K�>M�Q/�S_Z�	n�*h�2\.kaO���)�疺�㦃(�g�>���}A���b�%8hp�;���B���ߢ�`��9=�"�W�_�L�E��r���ϊ�p�fB�#�����9�.��ýSޚ�\Q��6�6�8�f���_�%e�,��^_��3�~�����ٽ�#-���{r�_�=iہ(/�b����1�VPȮ�W�;3�t�5�㖿�E��#G\�y^�2q�oŇM���٠�q���]T %*�~�_�fiߝJ^:�AҼ�kǗ�h�#j��#���~��<�2������O��qW޾�v@��R�#����� ����67�V���Bn��E�@9��;y�ջ��?�a����[w���-)A�4�V�lRD�vDr��,���Q9az�^9�$�z�y��S�����y�L�<�@,�g��(�i@)\H�0j��"��%�
1ê�V�K2���¡����-e�q	�&��\�mߺ⢶J7�����߄�J�Q ԗ0���	-���]$P5��g���w��. ��ʉz�.�\0��'ʅ���*-7��`��R��	F����<ZV)c�s:
�g�+4��/<
]Ҟ��R����r��(�N�4��x%0��i�$$�ÐVϠ�U�j���������e�=��~A/v,@�m~?�O�xgV��2��������$1�h��F�g��Yѻ����6������D���{�]��������iY��C�������rgS��y��W�^�������L��-�a�ϬWY��Y�-�v��ő^ɬY�E��ۛ����f�*�e�ⵝ�e�e��<kKV�n��Kii"���c�v5c�e'�ɨ��y������*g��x[d�s�W��Ocl|����&B�6k�ߺI�q�lV��m�q�d?��I�>b���Pq��u#G�e�.5Vr�1�{�ab$�}���
�~,��5������z����x��!X��fMlWMK!��oHP�~@�髊�-X-��yk_����� �Z�a��T:ɤ�n��D��-G8Fqu9� Jٓ"�T�%_�&{$�$n��̛�;cť
gS��17�2�b���B��:+�:�����s:t,�?�j��8�Mcni�sX��V g��2�*9�AO<�^�g�+s[�R<.�N�\�������Jg�%��B7���h�{5�6R3K��E�!�C��+p�,#�~��7�-ַ��y<^��,}|������ob��ɰ�_c��k�ߧ�_~t���,��q<���ڬ��w?�6�@��6�J�2�V�7� �R�D]�l~t�� ����>�x�zn��m�a�M���;Pa1t��U�=�uT��#�+����U�G��[)� $7j��೬�\�Ur@
M�Z�#�6Ĵ֫i��Yݿ9�Я��(�"%O���C�ؾb��8��JJ%f���K�跜��G���ҺG��
`GofF$_�ɉ|kÇ�����GםA�X&܎J�4�ie��aࢱE�oka\�����R���Xb�h����A}������)����Y�zC��zM����籮�f�M&>��q��A�&)���.eza3��C��8h��� t���������b��v�}�ޝ��O*^H���54T1i�w�����`��lA̤�S���!��1�_~K��dйP�8�ڸ~�f����|Uh
�<3�j0Sp��8p]�ث��k6�۝bR.޻���ɓ�t<��;�o��n_ۧA�*@��-A�_\�3��r�am���Y9el��y�|E�>�h���y ,��������N�������~z^k{)_Y,��I�(Ql�w�z}��
��n�e��b��]�p�rC�]|\"4��"�y��M������e!r����B�<������Z��e�����Q�ܚX�W�!Nr_��=F'�^d�ww��O؆�S~y��R�;l�8��2Њl�F6���)�ZPg���j'��`��vt5��vj�Sh v�7F��b�[�/hAJv��>:m���Gn����&D;K��<��#6�� 1q?���$���?�&4C����+fÒ&�O���wў������S��8n2�T�S����'�s�jqs��I�����6��,F���J6��m]Я��5��Q&�Zj��2�&E;���t�w{T7�� �}4�z�]쬛mWb\߅ ��;�� ���ٚ�?BD���S�斳�6O����>�H���-�{�����=�_�3��6S�kUg�u�X?�B�!M�
�L?G��B8����q=<T*!�s�,�������F�o�6l�od�<�4���m�*5�Rd����r�a��x����Re�1)*�D7�g#L���́���=�y��0�Ȁ����'��c�Qō�rH_U������s�S�%&3+<�7-ױ���A���Y�ž�`dQ�,��ܸjm�z��+�;�61����2�8J�0�<FR��w|Z���=��ZN"_�`S��G��ҡ-�����l���>s=�!�kڧMD��b�ERg)xE�|)�
y?{�;.�-��Gj��Mk'�2�U��4g�������7:�[��%EI��W0:�t�v���A	9��Z�ԍ�i��
{e�4�1᰸9!�g�h�<iǎ1�X0Do~�a��&���T�"ʀZf��=�qj�6nh�Q�J=;}�&�
?4�
.�]p���� ���d<bc���XGG}ˁ:T2$����
�N��*e|�'�-E�~`��?��@�aM�� 9�T��z�ѿ+*�	�Xg��l��R8��QPz��=*"C*�=Pp�PkwW҆�z���1x���8u^�'�ךӒ��)F�,x�$�|܆��� �l�O�8�:L�yM&�"J�X�אԜ�P���̌ ��.y܌3H=kE�iw�
{�Z9�Ԃغ�<0��C&@�9�����aJ����OT<V -,͎k���9eM�C\Ջ1 ��Ј���e�g��ŏ}�C0�;�4c�B���7`�l�زx���z\�wr����E]q쿮F�'�L
��ŎQ��Q�x	��Е[^����r�a�Nlr�U;(��6!�dl��y��:��Z�fN�GJ0ߍ����
.�갧p�3�b��SOLy����Bd�L�C.+��d��9�xr4%�r�C��X��l}e�m���!�.*;�����	$�y��k8��p++�h����$���{��|�O���?3X揁,�n��� ��Pݨ��j�lׄ:��#)�A���K�����׸����F�(Z��%���)Q��Hu<5Q��nEd�f�!��բH�A�m乩D�ӚB�WI�sY���ogeT�4���dv�d���!3>Zc$�{����P��l��rkOi�#׌}:�����a�u��+4��:�)��X�F*srRAW����fpz�6��n���fLɩ����s��o�x�x�܎1�u�|O�F�jxp��gL� ��o���	G*�B~��I�& $��w�mh�������b�����]0X琀���c=�	&�tP�<��$	�h[F��Q�0�&���uWW��"\ �rg���}�޶���Ğ�Jq�arͷ30u1_Ev��I����By/���;������Cƨ VS�����m�+v��-�}2��k��`E�٧��)���n"�#�߷}m�PX'K�o���]�?訟J8��wȶ/\��%��m-�T("bd=
��4WQ���e�1j�Mmc���U�qo���W�K4�b9��W]��1�m������gjư�|�n��]u��{y/�nxk��7�\�蟓�Ag�(~& 9 ���j3h���I���ȋҴ�LSe�Rs�χa)�Oy
�Ơ��\j�Q���@��n�_�	�aڏP��x>RHH�ȡ�ڇI��hm��[G�<��cm��ȧ=:��戦�p�� �&�ǲ7�K	aW~9@v�>�A����g�v�vK�v��	���x��r{]���*�5}��%���@0" ��_���Bh��k�M�s+��-�e
��g/�j$=mn6���J���Ƥ�XUf��������]��.,�Š0#æGE�֮���֓ܩ�-L ;K�C�<k2���\�.��u�2��:c��`}!��+�,�,�_�:_uv4�����<P�O���{�Z�Mt����'�8M���b�V�s O�-�j��.�����&����\�=�~Yr���b�&R���o��O0�5�ڶ���H��b�� ��g���<��7��a��5z�YpC_t>W����4�p,V��	8iB ����sY�����������h��x���,����k��١��-P�Y�*Ŷi{x7,����đᠸ�F�u�Wzr@��\]]�E2������9 �F]�&E1��눜��L�R"�7eE����.��p٨�>-���s3�p5f�І����t�n
��#�kFLzˬڙij4FHb�����3zFJ"����u�W�tݼ��֝Q,�ְ\(�����qۻ	�P��]:�,�?^�]��E���G\㐒���a� \�]�PhT�vWD@m���1O[7އʲ �|�w��6=~Q�j'���*����5���hԴ,�������d�j��uiV�K�sX�FH	5pX�K��*���	~^�� �o��q��]^u|ߡV� }/���O]��+2�*�d��p&z������ǒ�H���uMƹ0P���C(_eȆZ-I������ "C8��%�i���e����@�z��yJ������Fu��^�����Mu�,D=��܇5���˓�c�D�� ��w��f�}�Y����m`�e:+; l�yڹ4)�Pwj�n�H�]Q"6
��G����=lm�> ��Z�wH-SF"ֲ��$6N}�ty!~>bba&��5����闅�J)��i�K��}�t�����&m,�$P)6�B���ԙ�9Y-9�gS���Oy��Ķ¸|�^�̮N�`~���I�?���������BD(�� ������%�����(���]S.��7V~|� ��\w�f1	2�sۑrF����&g��zaa�%��"���/Z	�_��Ƃل��M�}���p�"���2Kx!�����b�=�ܚff�Nq�����^q㻈�u?��u�[5eg�['�!�$��Mu����!�y�G|k�;�W�;x���.��_Gc?�l8��HZ����A�*S�-�
Le%�wG,�o#>�FŦ���,��''���zb�/��,@�,_ćg݃v0	�y|0�F�L'�W�N���a�z5�b�S�������H�	-)���W�H�Pܙ /'�cOS#3��Gǂ�<l�JEŏ�����+!����/#JI�~q�f�ЀN��ب�H��Z�+�\�8�g3�q�#��̆�g%=x�vXs�)��~�����o�(�G�A�o���
�Y����ێ�K�TJ�)E�V̩���٥��Yg��Z	�{��>������VO����֏ycs�m�0~�ځ:�yЁs��I������~�~z2E��F�%��@���F���˻QT��(�Za�:Zɪ��> 
w���C���Im�����
봷��b�H�9��*���1�����8�5����`Xg��JH�k8(	�Ѫ����s�r�x����#盗���b���S�9)�@U7?�+��F����d�~�Z���oK^���5�G��F��-C��P5%z�fK�aa�Ϥ9<�n��� �����
�e����*'�E�7��-���n>���n����N����Q�0O��_4���H�O��%�׸�Ԯ!��s3�n�̀�7 ����0�;zK4��V�t�����BF܁�����	Iُ{�?�+�IjK|B�Ѓ�]'��)�B��K%�ӟ�*L���$Ȱ��؃Y8�E�Z�F�"�H8��$�b�w���g�
 p��/�ȌՄ�e҆�0�0��q{E��8��2& -r鰓�.�b�|~a�z�)S`� ��b2�à��n���5��R۪��i�?���M�V�y��y�H*=�?}�. �y����¡��V���;<�
��]0�6�?�c��؅��c��q�~gQ��̇�Nܿ��WMFy��s��cLy�s*K�V�ŷ�=}��D����t�?Eک�x��˚�.��.pZY��J[Pb>��ORn�T�]UW�AyB�o���Ц�Ƞ�i��dr��{F�ʠO��v�Ƹ�2�w�Gg�ϻ>�u��(!eet 9M��j�߳{��Ҡ�@n�r�1l<*���T]��+5�k��g�v��}c�k��2�1�(�dD�e��K��������{0K|�/�u���I�������Zm(��L!���M�h�QEp��:C��r�R�7J+\b�Lҍ�ӽ�xͥSd;x���_'�|_;jKo���1��#�ō򉇝�&;�]f��f?
��Q��>�;��+^��8^6�=_�ak2�FTqp����U�(���k�3^���%���&ͫ���`����ˣ�mr���<�`�w�s��}Hf�UE��/-Jؖ�{�p���guy��&1'+z�j�C��,bE�*?m:%�{�"����S%o�8����6���
H4%0�C@��"���Z��m������q����O �z1�fu̮��ᪿ���M��7�G�)0c�*ֶ˽�G��db����2rޟC��bY��
5�Ͱ氻\Tb��]{1e(l����0~���ϫ��G�w���a  L������pbh�aGG�e1Ʌ %�ȕ�vR��$@�5�Ի�����-����#�
ry\I����c��+^ƵO9 ��Yr9k�������KT�
j3��%z��h���6�#��?H|C��u)�h��`���p
�=V��&���N ���p��q�8}hn:Q�dM��M8�U�Y�*4���k�vp����&��W�u�!���=����������(臹S�q81��D5�И��p3Ě!�)�π"���Z���/��[�.Y������^o;����ϢG;���a��hp%<�3��t֢�h��%��|�c�º��^������Z��
_�����1�nA�b`kb�	���,��1�"]*XT�H6�1k����	H�,s���f��B�����J��]���~:%�h����vY�d��%8��ݧyƸ��Ӛ�~�U�u-��͙{pYo~����CQ�[+R)�e�+�tmR�\T^���ܩ6ٕ3��F�d8BF�~l~�G�(��^��ib�Hמ���� ��iY"
v8��f�)����Y�ږ-\��D��&�sn�̃/� D�>�!�b��C�s-�q��ڇB2��w��#A��A�7B ~~����5E4vh�r�L`A�Š%��D,����hJ�t坟�|]B�yx{����RԚPi5W-�u3Z�����`��ŋ���׬�|#*��s��g(9���|�sdmF�������<�Np;T�ɎLRu ��I�u@x������񽒯�c�WL$YE@"���?��<��G��z>���=6O6�8pDr�_����C��4pJ���[����@�	�2���nc�}V��"U\Q�m�[ke+k8WݝQ]	݆�7z�X�P1��T��p�M!�ə=��k�3/�eٜ*����u.�IIV���V�T�)��z��z��]x���\�L=P���p�N�w�K�w|�H� �r_.B��],���jm(2��^��q�P�%_�`j�r>o	yZf3�ddx���ݩ.12Y�y3�򙛭�R�g� AKՋ��e�7k�Ğ��Gh�XL�F*JC�Ϡ~~3J0���O��x�	�;�;��Ԓo�{E�[*ĮT4��]y����I�	�x����X���IQ8��@N�%/��'�����5�?@�T�^������Ir��؉[F�'��"P%�(4�Z�&�������3�fE�d�:� ^g�����'yэ䘞f:��WndZ��/%&9���0sɕy�n
(���f'��*oWb5�XC�I�l Z�g��L��h��}���Or��#N�d� )��6�U�����BQ5�X�QP���-:��!X%C��*��=�{��f���1����	"bp�oD���_��}�L�o |,)��a���h ��Q�5���܊3bƺ)�-��V�=��@/����q���i�1[41n`dk!TX�������I�qi{��	7>Ą%�i���7�y=�"-�+&/6=HYVԕ�)د�"��� �y���ݎ��C��o'�:�2������,�
�������r�;��q}l�}�ܖD�;5�8�p�l�X$yѱ咦�Z1���w���۴�j��KT�Rp�J������߇�,槂�� ��8�%�:Ƙ�&�9��3������'��MA
���*d�O� ԩ��@P�x��2�]׻p5���������J�]�Y�9����\����J��G��FLm� o�Y�HV���y�*�,�UM��g�D��2b��"�M�t��m��y��R����Y��Srv𠆍�/**D��[�/�Q
��Rkyv��P�����X�0�d&�z<��$&1k3&.=9�z\i�>�i:�=i_��R*���
-+W��Rm�F���t���Lu�Vn����*2�\n��0���q5��X�(�6]٬����_����D1DH�O�&ܤ����3z�|�řU���G��b�խ�E=i����r��lT��t������W�"�<Z:���"�Ξc�?-�x�Ѷ8\H�b�/.��)��w�k.x��W�9��}�9T3�6!�m��M-�7�"�T@P����~����������s�܋�#)�F�.�~�\H�2���4��<� ����!d�
���4�P��Ľ����ر�3�(�`�/��p��K � ?�!��e��{U�W������Q� �K��tw�i�c�IhfaEfR	P;i��8gc�	�e �q�c�`$����0�B�b�<��_d��:5���;* �Fi!>��]��K�C�f�k�|��e}\�'�6h!�uvcİdt��t�a�N:K�
�k�b#�G{�w����yO '|-�d�V�|)w�2(�R[Wc0Sj]�H+�ƫ��DΠ̷#�)I^�M����E�s��V5�v:�;�����Cy*o�W�����T��o᳟��w�1��,*R�_��7�W��n��9�]��4�-���F�$i�o�����YM�=����T��"�B�f�.��{!w��b���@%��9�N� �P�#�}�7/�X2Ӻ����H��;{�K�27#�6y	wt�����'�(n�;��%]���@�%�:�����/S�+[ɍ�K���i&ůs�UA�m���N��D�{�{���\����).�^9��f�|O-}WA4�w�_�R�����V��g�#��~ϛ�.�w�;�)���pU�:�Ӱ���9�vt���B���[������*��3��&=�QǗd�V���+l�6m�} U�>�lh�`��},��gȃ��S}`�_���xv1�J�Q�5'��W��*a{�M������\��9�n ���KM��l
\q&������f�¾�����W�c�\k۷̇]Z�-D#J�$�0�=��-h�C8x�����`�F���y����p�2�uq]'���^yH��ݣ�W��%���7��Gk}pRB\�X1��h��e�*����o1�t��Z9���P���Q�w�m#o��T����$&�d�BR��w���ክ�2��Sj�}�L.���C�~a�/�������3�ob��fH'�F�J�j�E	4W�VAC~J����vvw�HR����	��x�~R��ch���Se&qX�=��Ba�)��Mc7d��W�P-m2�]�Ո�($<l�	�Q}?[7�Q&FJ�<��цE�FO� ��Pe"�
+1��o� /I#�FH��O�$�9����4�� �^١־��C�O�yC����^)d�]�+�3[�Xs��`�o�Ņ�ؔ�5����T]����8�$V{*ޕ}��~GKxG
dND&�����WM�UNg`��*v�k�C�<���Vyf���U!)��/(�6��E 'R�c~Z2� �"�+�!��q�G���� 3�"s��s8}����������k�{&��0�!2;Շ�*��R0�� �bX��o$��,t�]dS�/lF1���+�E����*�O�xE��i����IZ�7�@���jd�E+��y{�./H�q��{��G�����]_�$�����1z2L�V�����W�I��*��yP/��Vg1-���^�5���������9� )�a��]*KEN���[ӂ�v#0s.�C6��4�f�D����y$��,����6
��K���i�v7��|�:^|I���ڋM�b��^��W ƚ�ht0����`N$t�"�.߫ZpB5�N��ԧm�V��$���xNg����l����j�I��4U���I���0ے���F�b_��Ð|���Y`��bf������X�e^�뾀jd0���2(�:�ڇ��3?U6���3���t|���?R(&�� ����r��V�]�ݛ�u�R�6��DZp��\��f�i��N�:�!�/.��5���d ωC�$�M-zX)�U�I�k��wx�vP�Xx�< �dW�xs�?�j),��6�?�eYNI�˼��in�fܭ�3�^�w�y��H0��Cxl�T�SϨ�kt.9�L3F�������!���7��b\���D�(�0EEe�nPSj�e��CI4Ѫg�;���T�Ρ�o��@��B��0�w��t4���S	S���Z��������:�s!=��_O���\���m�/�r��tGCfp��,�ל�b��zП<�(��z`���؞L`~�D~_���;�ܦ��$��\�ԕ)�-[G%��@3�2�b�/"����\��=cz�j���#�2Rf;� �N^/��\6)����T^~�4E�k���*��B��
	S�������W!����3���Ɨ1V�ֺI�jp:$�gj�� A? #�L�<=3�ދMY=�����EF9i��7��*)f�R�Sp*�7P$ �Em�$(WU�@Q�`�(h��I�+f����p����<�\�NG1�՜�V������������+���Z�_݂�m���g�_ZL%����<V7��iY.Sa�F 
��%2����%w�J�'����J��E����h���F]�����}�r��1ǽ_*0����^�3&�):�Z��t2�,�(6��'�J#ˡL_��g����iap���&���մ۷a�* ����Zq����]t���H=���ؙ��mM��=�������Z8Q:�B%��N��y o��.)c��oM)�S�f^���U���u������P�c�bO��G�N*��/r�)�-�I�LD:RQ����ܡE���s<�!}�k�,!���x�(UzxH;��XmX�$����?o��&��0e�H��P�އ�1�H,3�E���@�0|�^B;����V��\��:�:��&�AnO����Wݶr���/P�_ۡ�m]��O����@&���)
�S�N��P�"���9������t�y�M����>&Q��!9E�_��6F%2?9�P�����l��D>�ZK�4���z�f�}�a.��-U�[�!�r�d���N"�p?�;���X��!�Q�z��ri@p�*���#�Z�M��E�b/��wF\����� ��t�p�qL��V���qw��5���s_`6eF��p᳴�[�v�H����»8N���.�8�u�~�T�\2M���QlH6�Q�5x��N-�d��3tgK�e/���v�.d�y^�X���B��䩗z��X9���3���v[�}<�2I~l���|�(Pp:�p�bF$,�vȻ&���zL����XMj��+�m~��P{���X��l�v2�{o��4"�RZ'G�R&��������[�*�,�%�r�k�	�Q�p���Ҩ��dD^��q|4�#Om��R�D�-Ɖ�a���,��׶�;��M�{)rbN����tآ��`�3�!J\��Ӿc�j�?Z\�E-��5M�#H+~�7�y�����fշ���Q��_�m}팹��0�`�	+&�&Ү��`R������Gm�"Y�%F
r�����\����.�<Y��Tg�v��%�ɥ/�1��ؖ��*ƨ"ϕ�4 E�y{yĥ~�N���ŸMwG��@���L��\����=����޷��{���~_QJr���?���Z�u�� �a�Mf�OL`��VO� �@���D�j�/bQX��&!f���O;�P�Gg<��5~Φ;*��/�]���ȍ{��1�A��l�Fq+IZl�J���d�˛w8�#ޒi1hݍȨ\�����.jqCg�L:���%�Vd[2����5�О\�%���N��~9BcQ�������dV(nD���?%��0��>G�Ņk��m�|*��^Y��L���4
���ISw���j�|&����È+�G�䩯n��pԈL/q�HCJ�|{���)ŇR|?!f\ �[A3"i����k��Id^�n�x�y�ArD1bX����.�h$��X��Z��]%����6��xY����w2j� {��^� �?S�@�����А?�e��_��\�64H�RG�#�Q-in�3���qFlK:4h6�݄ko[�e �K���"'Y�df��� ���`7`Ml����(�{8�ᰙ���;9c�W5���nv����0�A
^�j����3\�5�5I����%!N�G�[b��Jܞ%�K����h��(�;*�高��+�� ���<�8n������ƙ�{��莈�°Ϧ���ϑ�Ro
*�X���R�Ä|������(������V�p�؟.��5�e9p�(rvL�I��F]zl�?t�e@�w4���]p�y��:W.@M��ͷ����
-��X��d��m@K�%I���[����n����3��� Xk]-��h�	�Q�
�>���0 ��cy����2|>�RĈDOM�Q�1�ڨ�1���X�^ܱu��昑�2͕_��t~��M�_S%��z�D���&���=�`jy�M�~7�[����c�MW7�vp��&w:s��|��ܪնt��O�Ubm��x�O���E����r[�`A����@�Ê��KN�ȑlf�:�%���t��י�^���"A�K$��L���r��"��}�)�҉��%���� d֑#�H�E���������A��ݟ��><�
���n���-���HR��=�nej�w$'��|��O��u=�F$�SX�2���"_�'�*Vpx9���g�fOO����$/&��E�~�PǶ1L�@&�u���4q��ޭ��)��m8g��%X 6���h�6�b]��ڃ���0)�l��}�"\)N2����DC`u��6�Vp�S�<+��I��]���o��@��kN��0���X-�"���İ=�Y�qܦ@ 8ᦔ��ž�z,oPx���X�L���Y���6��떞�ðt�������l2�9}霶h���U�� ������4�z�!�u�,�D�D�Q����]d&k�Y�W�Ţ���Q��b\��R9>y��ֽѩz�-$���(��\�V�(N�Q��(��W弞C!ܺ>���}	4���4�<�aD3��Yf�y=+ �ӄ����LA���>�J@ݗ���2���{�x�U��`�r��7[�Ff�c�Q�-O�A����O�3�o[% ����d$0룭�_�����m9v=�I���J�����w�'A�k�Y`�M�]�t6d_�����5i^���&�� �U����Fw�|9�{ĲA���~u�{ؖ��I�a��c�X�.$H�l��<�g��e)����9�����?d�58d8K�%�Y�˲�7�x��x����w�/afܖ�S�}��hTt.��`��叹]O�A P'\�ܵH�݅<}7�2���	c>������!��P�-�t��E׏K�A�=h2"��,�e"�ⱆ|���3���`>���8*�-��2wɘ]�I�'��vm�_̾|�F���zο�W�xS��u�¨�3�(D�:*~��EBJ�]��DWd��v.	�)�#ϛṄ!xD�_�����{^���Mk6��4A7%��wK��]�<ֽY�Q�lG	-��x�Vj��Yϖ�I��6�%Ef��M?�fğ$��%����4�?��Z��w������Yo�	̳� M����Ӏjx��m[]��F�gw TI�Ua-ӛ���׶��Tyg�C�a��0B�'g�+�F�XTo�XS$/�b��1�#����� :gl�t��9���v�D���d���]�*�^H�q�١ ���-%#�s��q���ޥ�­������g3�i�>@��JB��+_�rl�6o$s>;�����"�-T
[66B�E�&Q-c��՚Bo�.ɶ/`Ykr�{�zO0M�<�A��w����V��u��Ƹ��1RJ	(�4X���-�p�/�w1���箌A���-��R���Q_HH��P��bݓY3*Tظ��R)s��->Ce�#k�yz�o(8��� �W,�8�(���2������
@���~\�?����/����CО�UQr_Y;b���h�k���,��9^�]a���V�)pZ(��軹�^�w5�h�Q�T��:!� �ª���u�Y�U�nO7���ڬ٥���3}����Ƭ)��}ga��/�O��GYg�ڡ'����D�h)��VC.*�옔��m62`6���'��m��^�6Y߾�>���xo{�^f'զ˰:�j���%�Ю��̨1'�^ȼrU4� ��8�2f7�����W��y����B5���͋S��oh�-O��ڸk^�C���e��Ԇ��z�QJ"��}�[L���Q�C�~�(��Yjw+���D�ޙ��D��o&	 ���6�FA^��cLȚ�l�m?r�Y��EpO��3���˼aF=��H`a|G���u�IOB�~�K7T�L�A@�{e��wtz�?��5.�`/�4��V�)���^�4�щ���.�8��ܷ��� ؽ�L����Ls��x�G@���8���S��?����ATU����
@��� /�T�<�H���P��������T� ���"�����-a��C����8t!��ŵSEIfB�x_<���?�<[~}���f#����_-��Bn-��s/��_/�l��#��8X�Jp)��w�E�q�*��GR�K	q�s�Ҥ��L�-�E�`��	o-��bЕ���"��.�6^�I5-q΅y�/��&ي�d�Xl�s��#�qb>3��R3fg���R�7�xc����cľ� �3����Q�\��BqU���#1Dw��?���+�;�N:�K <���Y�/-�8>��VC)wx������n�VxWH7�j��x6U��P��]�G6��S,�|���p�6%a�`	�;�J��q
Jr�G�L�:�%v���h�.^KO��I0��_��p����}cGçW.dcM�N��'�ơf��և\Q�<��/�Ӏ�.��O�C/�f#�U\&P4:�@����-��*ńH��b�(����k��O��΁Y���{��8	�d)���Ho�;vw�����Й�ٱg�2W�;J �o�ɭ&�	!5Db�����N)�w�Q^� ?YL/���}Ud�*0��f�ǿ�}�ڿ?��Pү�M�|���I�7�wk"+T0]u����qvK��[$�Vw='�] �G�36r�~=��N��;�������%�J^��'��{�0�vf�|��ɭ���V C;��fjѥ;[I�8'ǋd�A#N]��)���F{Q|���؝M�M9��%������Ƭ�߮��{�uf�6�Q�7>���FDD�Pڔ(9�ʔ���Û�X�(#ҫ�"�c9@�y��q�ܬ�-��B�����:���Pc(�����J�I�,��^b/�����H��+p�4��h�#��ԩ/�l������K�>�j���4tU� �X��;�e�`��H��<�Xw#d��8�!���~%$0ۇ�����~���c!*�#3��&�oVF���S��cm���sy�f���قҪ��1tZC��}d�������#m"�JAoi��Bg�vt(Yx��Eյ�>l-�F�^r��rs�!S����&�C�Yy��� "Q%J�;�m'm��Ԅ��\yN>�`]$�MTp��Yțy�;�xߌ�2=� ,ٚ�蚋�zK%\ʊG^oN ~f_������c<X���{|��#������x�ږ>c �i�=��&B0��C#��Is�� 4�:�@:opv���"�?"�/�я �B��q�
t��
6	i&q5{>3��#��ö���`K��cR:�x0�l�r���)q��s:�P�����䑇L-��}��sR4mR<��L��s��}4|��+�d9?��r0�=��� ��x���,��w\�F���ʠE��HM�z�����59}�\3�G����I������2�(ר���c�������5~��=��Jk���쁁o�}I���8[		�/CM�C=�;�'ѿr�ڑ�b�]l�8-7�&9q%@�]�W��~%$ci�@�8�R&���%�]�Y����Ɲ���'c�q��':��LdC:�o����OC\�@���"mP������M;���'�̶ݬ\3>
���N��hw��0�:�c�tn����_�(a��0�oD�nhѩ
L�n@G�iώ���2�>Vr,�@���3���a��]T��"��ߊ]�<,V�7���~ ���"a���O��\����i�n��yjo(yM�ν�%���Ks\(����*?�Y��b��i�������H�c����j�LB������	��N4E���(:N�B������wN�8ts�i����] C������x���[����s(8f�|{b���hY��qz�}�J�ˡ����u�Hi4������cCя��,X�9�J!_H�;�CM�0��t�ۥ�I2�uH���������Mnb�E�[|�&�Y��y��DC�e<�mf��Y���	�����\T����ZQ!;����2p���N�@6���^�q=�&4��Ydî*3�!�;0Sh5����	z�YȧpNEq�h�<p��Q8���*~Dֆ���mw�yY�e�sAí{^'�!�+��T��ba�����Ee��8 o�0���LC�R��*5�������!<Fak����#��D>��ɀ�
�W��r�f��g���1��	�"�*:S�}b:���g���^�5_ez�e���B��u��_��Re��Y+t FT�R�	�,��o�_�N&k~p/p_%Ӆ��?2���-�-_�)
���J������R�6ڦ���&1��s-�ÿ�4�i��+72���2�X�q򋉜뚩gL��T��<��κ�d� ��5A���mg>�`L�(q;TE8Ӣ�BDIϽ�+�����U]�-~/H�w@���D澄����a�X�,#/��*�lNK���7�D]�Η
T��8b��Ѿ'Io�8�o�c��N2x����<�פ_�I�
w�s��f���-3��#��ћ��UZZ�+US�t�I�p�]�;��t)�Ɛ
�7��tղ�	�6��`61�=t�p���f�-ǃ�S�M��p�Q�՚)S�n�Cg������vz�������ۼ�!l����lD���Ьgͧ���j�O�ɨ2�ʾ��:`;�@��%sK�3D?ۤp��|2W{�Y�DP�y71��_��%`O���[�2C02�j	���We_�C�pcN�Y����o�V��-c��R��x�f限=��.�Q��{j MU,�(>��B�K	z:+��%K/�~�$M���z):���)��S�ʎƩ�V�(�;��mw�,���I��{����PK1�5t��Z��G��/R�v-�l�OL�aT͛<ĝ�ђ�Ҟ�i��PgS��,8[dQ<�IK�>��v]]i�'����`G����@�=r�w�.zZ���ڒE���6M����Pz?��aA�b���3�=�S�L]�0Ɨ�g����OV����ؿ��Bk��^ � ┸�߀�|Oz�S��ٹ&�a�MaI>�A'	Z~�����<�
�M�|(a�[�+�3���L���H�?>���琛N��v�ZA\��8�8��� �)$|t�}�8oA�,��4����?������䵍��dd�x�E�뇽�V�j�%���]��Y�����,×�R�b�g������Y�j�'V龎�� קZH�]%��b�Z�_�Qűd�?O��	���)F ��U^������K/�jz���ѭ�ߠ�]^1!��ﻘ���<�XjM��5̬��Q�!4�jXm0����7��DW�?<�N�x�C�s���_s*"W�E�!o�!@�z�}�F����P��	o�Y�u�HE�ǝ�z-����^k��t��d^?U�ƽڤ�*E6��!�$ܹ��@�0-������b���
���mbG���~�Z	ל����_���X��7vo���X6�$xc�׾�-�r�]6��Z�ÃW�䣂:��.��_�0�WVO�8`g�S\������/_������/W&ہh���*V�$�W�PY�9�ײ��Q���H��oB^�)�����zR��T�:"�^L�������������v��K�^o7��JO����mƬ��M8N�v��BO�V�j�����F�!^�q�e��hBv`�Mߢ�@�ܞ0b�켆ܣ�k!N1����e�}�#.9�Li-��u�"���q�L%�q�d�j[1-{ti�~+u:Y�qr�����L~C�T�l���]�;'>�M�hh�Xo_��L�G"lz�7�:-���JG1$V��"Y���?@�\�|4._�����3\�X�jz�z��-��d�}�#�L^σ�P3���ޢ��C�_2$ފ�

^����͸���&5�7Qk�F!��L5X�[F�iq�,�~��:&���E\�ju��1�Mly�5W�}�k�Ӻ�4���2Tl��[(�`s�(��K#`���Budy.k���h������x(|�<�^���d�m-ICY�T�f����T�b?�v�_iB�>�U.�qd��-Q�1w�^��O0|�p��_�>��a�y�����Xn�B|��3�*�Dpv���X�\��ٌǔ�u���2;��1��sFa7�e �x��c��?�cH����v���z�XA�U�0�ƨ�rml��ڢ��4[�$���z���x%�n��l�3�k�iz�c0�����������4�1U�5XДB\(~X�8��=��޲�@?B��9��a2��~1�_�f�#�=Y�N<dsI5:��;j�/������U�c��\�*�i�v-Vsp`ֹ�IE��;����0��بClW��Z\����"�$~�T@��S	@��/3�����k���j5�t���'W�]c�T[�wQ���'��W�	��w�3Sw������I!�	fqK�����<];�n��ÈN��� D���=�Ժ�o�ڪ1rQ�b�j|Z@��Q*�z:_�$\�n���rI�lq�[���h%�]q	�8܄���Q31����+�HnEG�Hu��l2!�2U�%͢d�\��!��Kax1[�@,~S���1��99k,݂/�4;���g	��jU��ҿG"�(���J��S̕�܅��k\�f��}�)XXzX�Q�A��͸��3LW�$ԫ<?�r$�m���867�߻ʉ�Q�im��g���l2�?��+����A/l�{)�ee�h�D�9_�x�8T�\F��5Su�Ю����]{��%�#tjo�~��-:ј������s^5�wK�c���]?Ț��O�\y�����s �w�V0?q�t�1%���n���2�`�ƨ�OЧ0\Qw(�]h�?K'\�Z��б\ڑ8_�:X�$�߰��{����j��
�&%�ǎ�|�*G^����!�=��Bp� �JQ�f&B�nwb@�>���a�!�EF�di\����/����\|�|��b��F�f�`礴��cI�=����0Zx�E��;�3���HL ��i�J�0(�5M��2�!Z��\�[,2�cj�������u���Y��0���'?�R�{#�}�a��.���ѓ�5�x7\D$�� ���k�ʈF5������e��$pt�4��A9np�1-��@��ad4����R�S� vL�&f��]K�߽`]2�{���5�X㵞�D��57o��C37���5K����E<ŕ�Ε�x�#�˗N_eP�&rYH����}<�4�n���©Ȃ
&��p�Ox�����Ȅ��V҂��R�?�z���	�3/�MdɈ���pZG��o����;У�V��ݏa��y
��� +�褭���4�;Hf>P����`�A��!Bʌ�}�^dg�.��Rq����	ӡ��O+Υ#m��t�L'��j��� ��gs9*1m��橿��V����!�U-w��g��B��=X��s{����7����\; 9U�5�˪�<�2D�W�#FOb�x{맪/{�ʇ}�ݢ��$�&����S�z�7�p*T�.�}�+��n���7i���0�KtT��>���I�1S���w��B$(�"d�,��d�)���\��nWB�ک�|�4ѱ@���aK���L���Fl@�h���=�����sO�ΦϭV*`�ԻY��3�h��`���`�����J�#��%*.ɨ�si`R���,��a�V�8�k�>�/���j��N�ǈxd�_�����3��z�J�*�Ȟ��Q���=��������vR�ؐ=��'IY�����j����7�6�l� T0��Wͣ��cD�``-sYX��/ު=x�"d�Xx��H�g9K�"��,{��=�  ��l@E�e��)�B����O���sZ��p��%Ʉ�<�a�<�9���z����Q�f#�O<�Y�\�&�d�}�>��YQ�כ����I��ڡ@b	�!l����	>��/,��p��^ȇ��O���a����-�o�I6�P�R^�blK�[�q�Hk�i���ׯ�.�W뱶]$�
�kW���I<�V��h�o�ي��P�M����uiй�➠��V���e~�	}����VoT({Or���������
�CyU�)�������V��A:�k�C.�D�u"���`#��p,��IQ�K�(F�>dbo�]Kgd��X���6J�o�#M���ן�mXS�ɝ�.Z"��\@KW�+/&H�	��Đ�&�=�&?��m_��Q��U^t+�
�e
�҃��pxY�l%T��6J,VEA��[]�);��4�T��Iy�ӕ���)2k
�Y� Ő���&i�cwg�u��W�t�I���2a��wX9
���m<� ��\�%7�p
�g5LȔ5o``�3���T��V*���%@a�<�!{`iSs��2�<!��Z��;�<I/��'�6�9������۲���/��t�S������*	��Q���!v��u�p���Q'�i��R�~�
V,�Q�Q||�!���AH�R�n �Q����'�L�c2!h�8T�?i�G��gq)t��ӧ\ "����:1�h��5��f��E�(�Ɣ	ζ��K�^Q�`����Vq�]\,�5�rSd����7�+�ֶ�I�xe���.0�\�z�;(�����2/q�.��d��q
'�	���犽���aTIp>/�^:�C�b��֫�UE�����	�ӳ��G=�#��#,=�D�t>�+O�q���h���c���޺�X���Gf��fvLh��g���W���9��O�m�H�������{G�l!u�w�TX�eڥ�����뫽���%�z��LH�	|�-"��B�Sh4 �(7%�q'��	p�L��?������Az(��ѩ�N��i�t��4�7^t>Q�p�e鏏{[��X��b���A�*џ�+5���ñ�Ta�gQ�`�����p�V<R��D\x�����d�+Y���0!%� ?��5���Y�~�.�Z��e���- ��S0iw�o�4�G��R��_����a�5�V��a�m�3�G�}!��M��/2s[������,�z��&܇�5c��¾��W{T>�(ۯA��M��7P�M��v�X�u,��k�����U���N�j���at�X�8T��j���e��u��HkqؾP�jI.I��5�&oj��خ�u���>H�T�Y�	��Ob�2B�Ֆ3d�E�{z�W�r���6��		���1�ao���l��ufM��7v�������Y�1�~_z�I,8j_UCo�8�Ĭ?B�K�i [��v��G�v��>W}�ݩ�+�A�sO���lu Q���%
hʎ�|}��+�����b8��?������J�eLh�Z=���[D��`�9��<x���7��j���sp�ė�mrhh~
C��<�����1���僳"��c^ Ʉ�	YZ*t0�Zo���3H��ҋcb�G4��}������F����8�.6ƲI�����
��A곔Ep������|������[1�v���3�r��|>Zj�)�	8�]m�]D�o����لN�z-����J�Dc/��ǚr@ԸJ�~���w����5ߔ=*�ts�ۥ��Yw�:�KV�1�ߝ�F1�:��Ve%�gXX����)b;\~w�$`��� �)��ᵽ�~�ǌWʋ|&�t��]���֔n;v[#]��r�-�Jy�଄��'�4~�v��%��)��������*p���U �ʺF�f�Kx������ ��I�]5_i��LV�	���YA8��T�̀�!�����jwryc�͑����h��=�������K�]˛-I�m�J���Ow_c�!������� �+W$��T��ܫ���<�|��P��gx�k�m��ާH��!��s;�t���Au��?(�ƞ{б�Ƿt���r	f��xI�K�v�AOУ���z� '����-�f�ǯ�ϴ�n�[��[=x2Q�8��tG�\}���,&J�o��(ǹ�{7�'���]V'��L q������G{~:8�^M�SP{<���%�9�g���z�&֐�o��g���H;�㤝�-�רh���⮑�Ͻ9�.�x�"���ίT�tJC���շ���n	���m���D/Dy+��.�)ʰ (��Z��(��k����3�r������p]&ܶ�7�7��쎹�b�{����Kq� �Z����ىr�[ՂZ9����sB����� �Q0��>��.��+�~��iSh/��W��@U�$R�:��5��$1����K�y�z�����LJ��?jI)�[n�Od�C��K��2�f�k��d
�m&� SLR�D8���5��)��g�hDn=���f/���I���d����:��Œ_52ܲ�+��Zaڱu ,E0�t��04���DZ�j�hN�ԁr�xOmvW��[w�5�f���+�i8X���k��K�s�sx�V"n����rr���9�u=Lx�V���r.��鲛�9��s�C�=�� �O,�p;IA��]y����F#�^��x�o�
Y0��*�!�E�AB���~����=J����!�{	 :-�@��b�F:�"�XF➼z��6cp(٩ ��b�V������Z@�sĶ9{Of�.W������jr��;Wc|p���:<�$��%��XSN�����Z�t�cl���3��Wjo�� ����uF��'u�6tQ���VO~?c���>�B�d)�2��j����_s,<6�e���o)�E��[�x�������
�A�H��gx�d�h>�Ã����ҷ�:*
��Yy�[)�5(�wBV��CS������_ W
fJ�;|��R�G ~�¢q�᷍B��N������IQ�Pg�[��3%�K)�@�O��7MRgorC�(���B�A`/�N�8D.�N с��"���� {�h7��,Gr��U���r�zEY+^�\yVҮ��r��[��[��Тl������b3c��X&�t�_~��bZ���j[H*95������EL�d]�HT*:ճ?
F�5�[�!~�8������+��A�zy���J�5is3"�:��3t7b�.<vr�K,�ެ�~}L02m�5��Tcn����}A~
����f��Nߌ���'��kڛ���H�v�p�+�
>T��%��7{�z)�ׂ��������{�S����T�)�{��4/m���'欋s_8���05蘞�P��)X=�5�X�����a��(o������Rl��$ys�z]Jr��k���Y�l��Ֆ�!ߡށ��|-�"cܗ �j՟h��U9tu'�7�<���R�gB���P�_w�|-ߛ�m�����}'����p0�|�������a�H9D4�>��+��zD�P&�?�
���3o���rB�v3�����OU|��?KG ��=�1������&g]W������������������9��"�r���h�����1Ȑ!��VHD��RG�����|=j-�?n��#J�g����d�� ?��W�U3�޼��$���}l����ԍ��Zj
���� ��\���%6X4�.)@۵����>"k٬O _sI6"z���(�oxAl�����rt���`Ţ꜡�'M��Wi�P��)ݔY�!�����S�ۅXh����I��$���3P�*�K�$��m����^5���f#�}�E��¢��; �k��q���F�I$�}��I�K�qL�=i+��p]e��P�E"��?���y��F#e�\v/ V�?Å�,ۤ��7X Ɣ	�J�ګ�t'm��6Is֤��>:��!�=�
Ҧ�5��&C|��N\ ��!,�1,h��~�E�s�$OSll��&E�'����`(�9�������(p���O'W/d���ʰ���$w���w�K�9�����'"������-��u��)H�P��I��s<�2/�Jw=� �O��e�AkX�V5�|��g?X�U�q\S�:��_Ë�_������i��7���UMzL�jUS̈	��WTBq�A1:L��{ k9���B#�-:o�+=,xP� �N9np.��A�����<��\LiyQq��e���<�ߝ��b����l�OMe�o�h:ݿr:���g�[/Rӧ��6�C1}�h�It�Kk8I���n[��;̳�0âViM8(����XD��Y P�X%��i��2���iG���-҂��f��������JP�9ũ�u��.���=̃B}n�x�OA�d�Od�9���OZ��=�����L�S��APYV��V��C.��jm�B����B�ג���jNr��MS�8k��J^c5�Z����ذ`�wBz#"o?H����b�ť�J\���,�����}��O�{58�����Y-ow�`�n[�m�g�x�FE)s�y����d����ӄ3|���c6|}�����o�(� �Z�zkc�Бl�n�&h��}GA�}�wkd+VԪ4IB�lw=��ZF��,uytf�9sK+���dΛ+�����r�7�x|�Q��E��fV0�H��ͺ@g�#�|M�$��t��
x���i���'��{�!8jAX_�!��Gӻn%��rx��Θ�G�����e��^�

Mr7|bWuͶ�X�xnq3���z�P<JL0�|0��man���b�Z��)�F�=��M�~-��'��~`k.z��bKU��JfE��K��e��SHJAI��J!�v���l�\׉v�6�ϚJ�E�+<��������wB	=�h��$:la��%D��Uķ~����F���4F���XԶ�1����nF(ZS����V�x��\^%�]��m�pߨ#�m
�4�͙}]�?����ٗ)�J"���O!y�]Ru������'��(��j��+]&8�k���U5�D� �`a��
n�Q��l�JZii
𼕛�b��t����c�N��\��gӟ����\����*���"��A�L�??{��^C\N��L�v�N������̠a���ڛ��7������p"w7z�O���� �����\��u�^V~">m
�|�l+1�6N�0�}cP��y!~T7Q��52ܬ����-�$�L����_�-�E�]�w���2�}$L͓��ݢ:����5\?��a�����l��t����KX�C��z�>g��\q�{�m�{ߡ��L���q����5�R��������H�� ���1����KR�c����@���f�t
1B���V^��!�R)�TZ=�k0N8  OO�ǎ�i�2�!��d���#q�v��@nӓ,
�\�$�U�WcA�I��Yb���7Wh���*'��~T�UV�t�A�f5�)D�/t�.o㭣���o y޵����4
�#�ى�� ��d2����Z�;�T�!�MB��O:�����>��������fŊt	�7�F-@���Rg����&X%|��x3�F��k�>V)�*:���A��ڌ}Yx[��H��Omǳ�'��'�:��S���:4�0xN�&��}�t�0O.�q Lb�E\�ֶ������M5N�����:� �ͱ6d�gy��'ב߃F����o�a�����F4�_���u�{�4�b�b �=��GMN)�/��݃�wi�݁�Xu�j���籆���j�?��Z��1�&�z��w�#����:��c�3�a	V}�T�$y�6���(
l���ms
U�gS��ߪ�3v�U7@��|D��Q���V����=��P�C�u�3,��Z��Dx��ׁXgk"u�-I���	K��n��B]��iD��S��s�n�_m��|
��@�Sس��Z�۝B�MaέM�O���S�_
��B\���\T�Qq7d�.��f}	`C�pB�Wi�4�B��9P��(�o���l�C�=�H�
�r&ќ�P�ĢGҎ��c��:���W�8գ �!p1g�~ai
�ʚI��/�Ja��J.���]1�i�Kq��"Y���2fV�ͻy
~���rn?�L��a9"@�O�4k�����H+yreH��3Q�v��s�G�j�� �u��K�l�Ǵ�X+��Qd��MK-�G���	��FGr�uf8�<(º�v��������4zØ���j��Xd��i38X2��w�'��_��z3��jɜ~���DD�в�@K]z�9��V��~�7�Ĭ%\'+|��y��%.�6���QE:Q��������;G��8EQ��`o���vd��-�(��q�����rp����J��.?�Gl�t���Z�'y�(+ɭ��WAӬ{��x�y�/�Y����¥���0������q��s�x�E8�G��H�T�
o��;��c��<�F�J��-�z}��M�|�0�֐qc�v��A��VHp�,h�!�@HP�������e�����E�;���z 6�M(I;�!߈, Ϧ[�q<��Μh���y��$�o���C�OK\#?iG��9��MwU�h�8@ꪝ�+m��{!p}Ϊ�fi����n-]7�c3���M�I�[ �A��j4W�<���s�B7If�ݭ�X���3�X ��M*WM��Q�]��XU�����1,�L�HQOny�vT�
Q�2B�w<O
�K��mJ@>e��-�]��I0?�B�a�!�I��7ǺY�/���t��ȼ�4a: �Gl��7a&�k�7$e�e;N��y&o3�%�|HUy���4�
�/�,m�'�)�5�d9���Ө&��"yB4�|Q����s������2nS�Hs
3��4�5i�{b_�	*�f�烤A�����yd-�tħ�r�X6l����&*c��@_�B���F�(��Rѳ��� ]��
r��b�Bg��K�-$��/�!�w{݃S�w8о݅�KR�,o���븖E����'o��"�o� L��N��$zx���ᣴ�t�L��o�T�Z�O�a�=i�qx)������>��&�tD�*��Եӿ�v�y.�n�l�Py`�<1ݕs���=u����z��*�DBp_q&��0���oa
0�$�@,���$P	����<�=)�m�42��V�ڍAbW%�S��s�\:��C?��L!���oG�Z#8Q����jYؚʾ�n� i�K��O����/�ʵ��H  �2$eo����K+�%�5`j�Y�n��K�'&�߄-P���6K�~�2"�dzq��Wt�؄-��9����rIhR9z$0�&�ƻl��`��4��B�bdNq�����ovh�_˧4֨l��u��)���o������X�H�4Em�W�4�a�m6-6v�˿�=y2�	?��zՙk��
{����TX��I\��s��B��N���S�7O	{Ɓ;DD�M2Y��ޮX�	��QQ�c�W���,�{������if�%TLL\:J�Ҡʭ�tSi�}����;�����@U�
�_�)�É=���ծ�w�6���EqW��1������1V1c�#\m��0C	wt'F=bh�D���Ú�f�\҃<��e�ɪTU�}���1.���!{�=�Ɨ��f|�.�����0��|_�S�E�c9/e����q��J��j���܄�L[�쿮���}'�2:�J�Z����E�O��a
��V��^O��9e�hy�F�ga���ECh}�xWK�&�d�hy�+^��$�d������^�B��I��,�\U��,��v�Cռȧ;Vʤ��x�|r��>�\����=�<UԂke|�֍�@���:�$��Z?�P�n�6Z�wn,E���Öq����e���a&_	�}�r����#8�l~�K���`%J)U����[`��H��!mܤ�Qڐ�������jj")��e�Z�*�EʎR�s%����~S�_'�ō��!I�͍�L\��c���*���$��1?��q�E�ϢɞҤ+(�&�V/8<L��Ud��Һ���V.����a���}�	�g!���pwZ)�O�XDgA�+D����#�%$��=�}`�lV�����8W����)A"��`�>6?�#����~0o��Bp��$槳�>q�L�o\�(�#q;��I\��KY�i����D�Π��</��ўr!I��������|B����Mr�,�IK�jvl�����Oe
I4
�t0^��m��������,)��w|���<d8f1��Ѹ�@�7Xr<:��?!|�PF� �w���7
�c�K6��@��i!��'��h18����м�q�M[�(����]#o`���"�oAVrW����!q.���eq����b��M�U��l�"waǈ���� ��s6g_�����J�xu?F O�y)�׬�)	��k#�.m���04�� *��R#��<��C�=4���%�+2&]��y���BgDy@�O��o�6��s�g��7N�'ۜ�������}����kN�g҆����QxZ�g��Ъ��|�/:?5L������NC�{(��QR!���"��OT�B��u�����(ta=���l���o].��]̹�Y�__�Kg��?��@"C�7�,y�k�KO�N���޵0�m�F�O��r-��1���<^')�v�V��eA�8�~�4^dG1����uF�\1�P��7Q#�i�]85We]���V	�j&�l_Nxf����<��%�צ�D#��6Cv��r A!֓��c���W�L�쩰,�aS#ضdۨUص�-��%�Uؾ4
�"��� Y�8��·�**{A��K�g�T��B��_���,���[�����d�q�J�>	{/</�1�X~���E��gxc��m�d�~��7o�	���e��%�,a>Qn�@% _,�n	�Mw����/����T����#�i;�>0j��(l��Ia~`<e71�
>�E+C�� �z46�?�����KI	��n6�I,�䆝Qf�T��_1��G���
�\�DC̆&�JQ�-�'�@��/�'��%�~�e(2�[():j�������)ɿ�v\#N�S�M/���K������x�����\� ���i����º@��4LS	�X�K��X	�>e�y�:�ϯT,q-�Ӂ>�~�-i��``<��yh�*�U�GX	2h̀�Fy�
OsV&U����w_-�P��ui/�r�cVobn�V���:~M��"�ޏ� �Pl�]}6���a�ei0��sᾍU���!�,��cE���
�& �u��޽B��C�)L��>��X"�t޸\�\u�����ט��b�1�>��
�� ر��_�D�3�pG�<�o�Ǣ+@��[98j�[F��#�L���|���(�v�?��HF��-��f`�e9���b ��u��O��[���EeP�+�}Ƽ?A��(1˳�y��`��g+E�<V_$��^��}9�\��8�"�c�T��g��w��)Jw�����Q�V� ���B"�)�N*KD)�{t�V�Z(z}��i��4��C���<�6]v�ꁠq�̥(�V���
�׷n�w�9/�c��uz�,��ݒ��f�����bsq��������UkI�iR !�(N�@�/��K-�0V�,oc�W����ո/�7�d�*1-��[IR� �W_,�j����������eX�r5��8�'���O����p��(ڰ�P)��A���nN�Ii�ez\]v� ��d8�T��K�YU��kZ�y�D��Q��BB�w����G����\87%�vE?��x�ttvk�ϐ(K}�*u��s�����������mS�$'��"js�+`�6�f|���hhtH%�"�`+�L��
�j�>Aq�a��,w��;ί�
��Ʋ�H�[�Q��\���ᣅ�W�n���r(�)��X�kmG9�^�.iN\�7!��Pg��Nl6Dƿ����S���?��Wl*(p0lА������JQ���&L=����<���K�J��w��#�|3eWT�<V䵼BdYYq$�i4��ذ�W�'��s�	�����Hc�n��y���l �>9B6�J��@���ֶA����w[s�K���4֓�;o\��VUy��g�J�<�JQČ����,�K�ߤA��t	�G���r��K��Y���0�%4����[� �1f����R"0�.Q�dV)��|�?����"0'�)F�I�-�J�Ah���g]o>
��?b��mQƈ�����z^������1̿��M�d����.u�_
[]T��Y juh6:E�7'}Q)d��T��ces�I
�+~��pЧ'�?��h����|8=;~cĲ�[{��'H�y|҃�jgf�0�G�2D�8�M��AA�b���6_)Bl�U^3�d�K��޿��:�}��G4�	7��$Zq����͝L�ɦGPN��H >�ÿ����&\�E�޼�y�Wg��0���\do/����{�4�G�'6�`R��&�Y����0��@��O�_�=��	�Y�J��޼��<8�)�=�|�2��*T����G�g�� "����M��ܿ^2��o�+����.��f����]G����֮2��F���T��A��)�ܡ��vn���o#�f�@�53�Q�ԣ?Z*���sr���P��p�����<�튽��&�k�CKT,��#��7_s�D��'��텔n�2�T�X{�H�byI��f��
����J����������rsM�@��|s��f5h���J/7�J�&2<�ިN��Fr�<�=��;1c9h��,�zB	��).s��ԡ%�U�L����C��l�a ��Cu\�@�������y��M���
��@4�r��W!X�v>^S�kf��e �{��]�ep̺1�S0�S7��>�D��J{sE8��k3�§hb�Ɂ�.F��:�?�	歺}@�ť��+���v]���`9���Ua��͌3�������a��a|��}��꒦�ѓG�,�i�����2nd�ݮ�PN�Q%��Vܤ�SiN	)��q	��HujQ�'���:�Nly�e&�k��/}B%�� �x��4W�sV牀"����栚��"�k�E~�j�z�����/&}"�N��J0T�ԗ����(�C�#YF.r�|��o�$"6v�=0�C(HoR ����Z([V�}�@Z����ш$5�MZtq@x�ȩ��;8N���Z�9���|d!��W;��wL�M�� bb�P�6�\�=0>�ޭW�9�B�%<�J���
��i���\�xb�-A�(� �%��l����V�ʄ��¿䴇_	;6�!!2�eiȲ~�5���Eu_�]���S��{��IW��y����y�il��]�����*J�U�D�����D�T�-zh�㌼,�a�����Rf���]pv�#��*0抵b�}CM���"+Ϩ0��l��*pb�Y�M/��k��d:HK�$}rQmZ��x�s�1C���� z	4q���Qq�cH#M'�E�<H����׷t���p>aؓ�د_�Pb��w�D��78�y��2��v����ֻ)�
��Z�����	��J3����7h��#���	���j!I/|�V#힅��|�=�e�<��U���0Hj��U��B���C�<Z���I������7:$�]~]���´�Z��K��)J'��	�d�W�O��\O� ���gǆPR|?xړ�zk3/[t7ؕ�Ԅ�|S�(��Kq���;ZM
+�8���'-�_�55��umx���g��q�\`��%�w��������$]�L�,����Zl�TU����������q�˜)8QP��K������M�ރ�j��0��0z˾"��Y��\���`:�����l������AcQcT0�̇A�Ddb9�}��M�`{�X������ϓ�����W&�]��m}�p.�:�:C݂f���tbL4���T'q-�y��A��bH��+���g�2�������@F��P�"�qt!��/Ϩi;�&����VQ?��t����釥#'r+"�D)0�NFw�m����Q��p4;�5\����]V;��f�)����k�Hu�	xS��'��Ta|�I9V�N>5��;e�ӓ}xC�c��^#b֕XX*q��GɄ�Uc��%�g��AfF(�����wW:$m�Ƞ&ʪ<��$�G�����*u�Ԁ�1/��1��pd�ed����rU��.�A"I�Fd��WW���G�^n�b7D�Ǖt�j|�2dJR�Y��N��Y�ƫ�&��ǟm"��H9�׵�-Jޮ�[��$ P �+&4a��|o��?��Ne�!��z�)�Po[�	"���U��5�U��M�o�t������<�͝��d��Cp_S�m���V3wǇ�f�m�����L3Ԝ�����Vsv/e�����L����R�<���b�2�9��#?77��2u����rF����q��h7�q�1��Ƶ�x��D���89wѤ)>O���~��b����cw�v4��&S1ӂ��ó�r��h�\�C�|w�(��a}��N�8�4%��8o���6�b.����,���`>���״,�[�6>��oP�W$ TD���p��K�)j{3X����HP09����۶��OM����+�w��+���9u�ve$N[/��it��e�i�[�R��:<����6�!�c��>S��E�C.�|"�y2\�:�'u��tUH�)�[CU
�E���h~�3�3�"��`<���6�؋�ZU%�����Kd6�� �#�̾g��9��	�H��=Sg�Q�B^�Z��.S-�$�����$FE��Udq�s*	 ����ˁ�^�O�S��dtȢ�N�����Qr�oy��C(ř�W0�R�-��,�'����>�����ګ�1���/�����X/9z�
Ի$*���'QN�(�lS��F���r�i�Y!Z1�Y�����u����E%l��6��IS�׷h����Z�3�W>��z�9}ڨ�k�P��z���ܷMQ�A���r��<�c<Ǧ�o�mHSOv�s{M,юp�S?7qF�``l�H[U8\�\��\.�'��)��$�A߻8��Z��=���L��Xυ���L?0��r�蹰L����z���Ϋ���q�i!��Z��)�� *uUmʁЉʤ��t����!Y7�������%U5�'O2��~ܐ��v3��ʍ��b����~\v�kɵ2�c���Է�垊���H�*L��'Oq<�8Uf��${���}��KV���S]!|Z:�{�8�x�S��Ƌ��˯�K��Q��׺Fݿ5$���d&��`���M��Ld�O�x"�)���ƴ�BA5���^ ����|�L���O��I��!��THx��B��O-�S�Pφ%&~l7��;Z�t~�?ޥLEJ�<�Z�kE���v�j��G��
��l�����]&�7(7:�sC����IxITdD���W�?�Sx�%R}ڗ�o�*m��5#�l���WVQE-��F��l$0v��i��������/�v�%�`ox�*+��V5�	J�>tP�X���{�s���p��
]�#�w���p4����TT��g��g��K����s�h,xMGEw��	j�_C��&ȵ�7�y��|[�"*�׉}���S񟊐���E|�k���mLi�YPH���ˌv:=��I���caT�%�+q���![F~!Y���v�g<S'k�qő�7}Ӊy�l��4G��:nkp���5f�_�S��)�?B١�ɞ�gvҭ^�<i�@��W��7nna���e"��*��jۏ<D`mЛ�_G���.c�������^,f��>9���jsq�R<�б�'�dB1?��wCۚ��F�RT֒^Ӊ_1�+��f%L����7�����wa�
^�Gz�=&q3.�|$aQ���@b�ݔ�z!�P7^��a��hu��n�X�+��c������q����M����݂�77�#]���)��#�h�2��w��we\�����1�Ϻ��.q��Y��<K�f�C�6�ӷ��taU����,��y���ݖM�Y:����0��D���Y �&�3�Ƒ�V(s�DQ^�G'(u���B��,���z�O�&%�x?@�nn��=~�ë���5P�:<�%J��u�o�X�5~t1K��rX��X�7�zqR����I����ɩR/T6�àS�M�gX�}����/x�ь��5�+<N��Ĳ(1B�����aAء�c�C�b0S(��kp�ș�M[�����������n5�'��{��#���x3�4FW�5�żq�9�������9�t�.)�y��G�4��+�)����\5��ꟻ't�)u�5T�vU��N�<�
gE����~�O�vS��7o������o���+0�Nb�qM�F�@�`��?63�Nl$/�I�%27�����ξ�P���[h�:��dQb1��X�lZ�K3f��=�텬"��^�3N���:����l�f������<.x��X�n�����є�t ��o]j#D�:'c��7��ږ�W6�,�xY*�@�vLQ�a%�SC�,���p�dB9��2�_ym��.4w�y�V��g�1��6񦄳S�0+X���j[��T�U8���Ċ�s��<���-���+@ux�,@���9�J��E�y���}/�"�I$͊+켫��%�]�����;S`X�h&w�aUҒ2�{�R,�bb�@�eo�!k>u`Ux�v�-b;�3�����-BA/�P�z�x�����%�?��sI�%��03�)zL��^�
���)Y�F� ʙʙ��.���h�Y�AI{,cL�)6�T��Kv�W��RW�� x~�Sm�W�F#�|��@Tg���P�מj�ږ��*��'��p��su���uYх�@���b���I�AF�ϙ担+Ww|�A�z8}I=g�`��lq�ė�#{n�ݤ�"7b
�ί����06��� 4�O�0��̆~��e��hs�u��N�kV}:i��[�1ZD�"
�F�Z�"�Z'��f�d�[��W�i�����C�Y���Z�A#��/G��G�3'��_9�aw�O�%�&6B��5�d�&a�k����lXl���4��@n��$�_x<��vf̿�"w�������J�	�g�����(��܇-�����v���a��PD,1�<#�^����%ŕ]�����ܷ��ņ2~:]���������l��%vak��R�<�l�|H�����i�C/Z�:6���$�z����z�jom�H���f���&pSe�}Ҕ��e̽R@ �$�l��<T#�-oTl/�=f�-���<������5��O�ΊǍ���C��Rk��.\�~�����F'S+�Gn���!��sWfg1�^|�T7Mj.�����`Ȟ�3�ڙ�"Z�LN�L�t
,�kv�fU��K�JR&	�8���Q\T������v�Bg��x��e�?|;����=�s vX)΄��'s��Kv�rݑ��j��[I�8���v4����WQ�l���W�̿�4��%�c[�]�57b�"i�9q��N��uF�:�����n-Ei}�p�䐺���]Ħbl?�<I�`'��2���A>�w�����M��=z>��SX&o)p�5?��ᾒrO����ש�d������:D�s4��.cx8�7�s�>,<w2S���a�tƸ��I��[�<��t�8��{��8�3����+����D2�(b!!jU��w�Ѡj��uv
Q��g����G���A�Z���+��d��O7iX�5��`gAG�ą�M�`�{���u��43>�%߾��}ɶ��-qR�&;����6Xd�3�D.r��a>�a��w�|�x���d��pN�ͥ�I�F������֮�A��F�v0�r4�43��q˄�E0��R���� �Ҡ'ޠq}h-��C�~�&�f6h�}����('���ԁKL�Ժ�	��&K]*�)%N��)ɞ��ܻ��KV�8�r�&�,��фz?���$1Nu_g��zһ g�Up�)7d3)j�)�dh���J��L���?�k�c����]c��r�u�,��/A#n3ݢ.t�����{M��I�f��Ӽ���/� 4�{�h��:�A��D5p���~�,Ht�\��4�&Vp'Ӏb���?��7cDW�쓎�:��L��[Q�_(�9�U��^�^����%����]
��5[���/�� ���ڟf��r���<�{��o[$%^w�H�]k������ϥ�l����c9d=��Ň6L�9F��v3��VSo�I���m,���%�z�����w�L�"�3z� 0��.�w\��x�$�xU|WN��s�JP�a��|G�,�N��ط��r��!6�c1g�[�}�_�S�f�<��β�5��^�I�;�����l���?�S.�XgN��+^g�/��D�����V�**j+vǽ������Y�g�N���:��0�qO�B��W���1Ȁd�����K\��5����w�/��;�����a���2$��ڑ���jfc��+��p�B��拿$F�AK�6ͤ^m�x�f�h.��4l�hR�5y�E�wT#��&��v�R���m�\>�W@�j}cU4��oB��ƭ�i���e!�*�,Cu���jdr�~��ZQ������#�D(	��#)��p9SU8���W�C�~���TT�����f�џ5�x.�x�q.K�4�:�Һ/���H�&��7���P�р~ڹ���d��bם�T�k�S��'��c<R���?sk����j��~�����見!E��(�PT�l��"�� � C��R�&�˘��K�<�r|ڒ����O/O�2+�aLL���Ɲ��)�A�i���շŤ%AT&������;ލ���
/��9:�+�a*�3�@'��04 �xY<���+�k`��7^���?ⵢVu_/�c@��5���<��6P�~l���N����7���BW-�4;�>��4�%�\x�zaOla'�0�P܅$-i��>�d�3�ZbtD�w���j�s�x��,Ej^����|��]Q-yd~�.6D����aeơ��ɺ�0����
��M�n�!�1�����R/���t�N"�e:�����=��7����t�8I���ìJ��T��Zw0f�	�h����f!�9�b�g �ɝhڡ���ܻ`|�M0�� �J@���*O,��Mb��d4TK��<P�ow�
/�|v��?F�֛�h��R��t���Bi�Ki�Ԑ`�}���-��EGN��!R\3yV�1.���yZy�� '��:�
4�&�F0u���2D?D���RD���~�{�P�m[M�@UH�[�X̦��}�v�&= �<x���[]�l��Y�㳣ı{`��R�r�vx�ߍ�)�7!y����	��-��1�%7Ӎ�1Ħ����m5Iˉ���2c]ݦ�|�~H��^�j�_����^Me]��S��U�G�X�1eh����J���WFU�=E�����Fh4��D�]��
��{J߳�ҏ/�����i�@�s���$آ��u{�����Ȁ$@�K��A=FƄ�$�!�����]��#�A�F@��҆�(M�0��	�U ԏ��:J�(�=.����mM��dXf�(0̖?O>;礪���#�=2�B�X|g�i��@�%�Pg���B��c��)eز|S�i]�v��i����'>�Д6�S��9Q��C�}�j�c}~ףg`A�+̆"br�P1�XǢ!�O�0M�� UhQ�-����4�e�q�a[���pdM���h��U�C� �qT\p�l�ڞ+n�GzCpʪ.��*��eR$/~D�Z�ޝѯ��UT
D��CZ=1�n�0��T�sW�����p��x�5J��-fjC�(����W�?D�>�'㬃j�Ieul�ĩ�T$X�)}���,���Xb�3��R��͢AO�b�J����;�Y�~gJ�3s΄���e�K�/������8+���@�{ �8:�x@�?/���2������)Z$#I�8��W��)+j�Z#��8���W� RI�!r4��hv.�9K�8�(D�6���5��K$��t�O��N������Ȥw��nxl�&)>�+��~$�e�B���x؄����o:t��u|?B�^���/���K{ix��Q���פ��v�L`�B_��[�R5�2��� ��-�t�i����]ҲjT��ID�h�l�Ӳ]�b�V��	�'�Kר��k�\�3c���%h@�E����w�!*C:Pt�DO#��1����I:����U!��1���RM���-�Pw���Nc��f�t��F\���Ho��}����m��a��|&���J)D~	�m`v��%,�+��#��F	����H��0 ��{9jnS�5�s��m>*]��ꁏ%�{�Mg%������ݐ	��.D�
�?Ѱ�� E߈]5�p���1�D�m�
2�[��"Ģ�f��=�����F�B��I�ޤ%�����^���d�ׅf�\�z�Y�a�|6�
�����dezPd���&�4�/4�;��S7{8]��Gi�h��*F����D�M�w���"?0�TOJ<$m�oj�eV�G�|�0���vLѠ1���� �0��p��%�F��$s|�������%Ug����Y��J��RƝV�z��֖�A`jF�a��zMx?�@�Y���Q�C̚d)+n��RR���ڻaw�5���E{:��%�u8[c%�vTn�B�C�ܞ��
<��
�J�#�Ą�N�!�U�bw$��ҵ)l�6r`t�W�@6@����a{d,�B+84-?��
��� ��pZ9ʍB��~ 2/]���\��]~�Q��|���'�(OQ`�Q��F���q�E!1�C7�hvC���j�c{$���U��+W�o5^�v�al�	to�)�裷�!�>��k�H��]�"�hA������F���EF��z��85��M��Moc٭�����[₏�w>�y9o)q����M��Mm�h����=�w]�4}�ˡz����3��3���Ҷ|��y�aа�K�Ee)�6��[3�����3��ڱIR_Yڵn���G9����p_�^W445]E����H�D'�hp�a6u���~�n"u�T�q12T��l!+ʽ����d�?]���Fx�0�Z ����^E��*V�߽n�q	�b-���+W����[]s&j��	�j.V�ҟ�$&@ys֎Yi��!���C�wq��V�&[>���LI��ǉ%�:��A�Ҧ�+�{��q:�x*	2��_&������4�ȟI��7�pWiX�����,�B9M�����Z��凪fU+/����k)�
	\�� �a����w@I���#k�|OVL��?�CY��Q||���	���6#Z+�b�0�X�^����)�lI@���f����,����g�U���k)�d{�U��.�߇Cgw�
�V���{lZSԻTK6��-�&#/T�;1AP���;]��cj}o�� �j:�/5g�*`U��h�{�N���-'��,�}qb�B���?Ie~�FXL3���l��[a����d]#C��������/�<kc�p����2C�C@њ������Q��
޶�����ӏZR�8_��!���ѧ�D�o��m�w��L��"��"t���[��v�.�qy�	�@�XLN�,�%*гuS�D�)�|��'��_�7�E�Ӯ:2^+ �6����k���
��]�s���~�l7��X��/=�D���Bu�j��P��P+�G�w�"%�gcvX0OtZ�;�t2(y��tG�-͏��3�;�����R!M��i�Q���*T�ɽ�/@�����{��< a1�.gM.�'�M��� f"�7<�AI�-�w�����:�;RZ
{���\q��[������<�rD1���K$V&��S������Պfݍ[l(��ͧ�KEO\y_底fKQv&���;�ii"!���$������}�[�2����6z�jIx�:0
|�M��^��2;����(��쮞��K�}3y�>;�T�����w��is^a�/��8�a?tA��y����Nۡ_�p��.�6���RMݷ4Z���~]U���;�]�A!�����U�y�����z%t3lR4sG��Rec0��S�Ԭ�Z����c�����uXO�z(݇�-DoRh{e�Q����9�X�8Y���썮zՓ o����E�y�= �@4#�O�	/��c]z��Px�:D����X#�"&�7!=;���i}��
��L���4_V�w�9��JZtJ�EkM�̝tM;��=���|,5E�l}W���W�.�����MK#�M���P�[V����h�2�^#���3��|�����3�<�|��jt��]�Ԓ�zV9�'WC����'6�u	<\~e**pcy+������Φ�%�$�3N�7���P� .y� ��H5J"��8R�|9r�
6P3m���!�}�����.ÁR�	~��L���3�r*$��N ��Za�c�ab!Pay���� �����DW`�A�����x�Q<x�k�E�XX�	�t����M�3ؽ��]���m{�������NB��Nb��� b�QC�Gs����ķ�F"O����x-�� ���QA��H;96�8��;�}\�,���q��S*�kX}�0+\����q)��̭t�=7v&��2}�[�L�������'�D��Ԍ:���hq�L`�ԟ�e-˭�l��_� ��4Y�l�V��[��uC�<��B��X�H�E�z�9Q�Pқ̆^�����V~��;�� g������0d
��>�<�[$a��hW ���d������=�{>k�Qs��ǘ��`#��(��Y h=��K��:�(G#(֚se���$I�ih䙤��p`�N�O��j�i��R�-���PR-:{��)J)����ݰ0�	=���d�S�+��ڶD�#'5��/����%� ���Ȉ�,�@<����xї�I�h���g�xϹW?#�N{F��	7�A��	C1,�Z*�y��A�t��z��A0���/y�|��|/��ji�c��㓙��.��Sя\�~����b !�R,�E+�	f��:O�YTT�/|�R�LS�إNG�Ft���c�I���N�m�j���4�A'�-���X.�X=�t{3�m����n�3f��8ŉ�i��_�)XD�n�;���P�[��FX�(X���x���o^�	v#�3�y��9Xa�!	t�݄�G�"�=X���\Kq�����V~[��.]»)2q�;��b`V��ga�,;M��!�F(��t����f>�G�K�C	?���Il;�����t�u̴/�Xb�����TM�[k��(����>����(� cg��BN�]�4���Z��lS�A�/ޚ��Đ�}O���BV��}�h�y,���]�����I��$a����Ǌ�Cu$`M
=kgw?ױ�����_���Α�~B���/�}��}�D߲2��2�an����8e�i��E�؟��x	�$_p/!L���"=��G�י�;���S�ߝ.5r�^�1�1�~�EP�mQ#謺�;x�F�y5f}����� gyԨg��*s�>T��dĎ���	ą��j����i:rϱdF���Uş���%[��*K2eG{�Z�<���_�
ԅG�� �������Wz~;]�#TA�W�r��[�u��[�{�!�Y[�y?>lהdzV���rձ*&��Ղ�"�$���=%3���X]11t�w�в��9ϒ/G�9�͝��З�AЙ��6Lp)lX�Uv��2<��e�Bxt�~��%Wi�R�����^g�c/�� a��������y?o ɽR���>��G�=�8:x�`-u�A�̔�[fuQ�ǣ3�mj�)��/rĸ+>}D��t'�؆�V�!�IX�8ꄁ�?>��	�]S� �T	����5ߘ1���N1�C���>��i���[��@j|�<Z�@��:!�C���=Oq��1Y�06�҈��D]�1���!M^c�"�� �+�>��r�T=,8������e��4S�챣�ΤiEܟ�m�y�c^r�c��?TA�d�;YWZ��۔�A�ר
|�Q��]Z5�Yw���Ei����F���s�1��:�a���&T���Њ���^\��s�yd.��Ԑ�g����>�Lㆵ!L�w�dB�Ŕ�#@��ﺨ��vuɧ��,������_�3����` �&N}>��k�����l�x�X}�p��1�Ά�o���2��=ѥ��w3�S7+˹�P�Kc��č�bÁ���]e��ޥ�����m�����n��CҦ�)�=�E�ݢ�Cb��_/�.��{N��[�.�v�a!ZF�a�U�Нy��{P��A��Q0�v�
�%�];�<aG�%G{���:��`6���r��㏭+��t��+���ڕ�����MRq�����}D��Ǩ��{�*�	Y�8p!hh얏hl��qF��>^n
:w˩Z�s�a��d� ���� ���*�!V�[��T�u����f���]�l��7��T�-��BVktQ f�W�����Fj���B#�>���5�r`��e�W]��
�}�� �M6�Cu'q<[l_D_��Z��0�f(LF��7!��Udy��6 I@�N�ax��`Uք��o��r˼9(hM6x#��&���K�_I���nxZ4]+lIRi$~D�\�8[~�j��luz?�Cw���[m�hȲO����τ�A�Di�40]�qJ�}�i:p�uuf�A��9X/���$��r�җJ�:�,�4ad��J�Oo����D��l���� �3�C�-��͌�������H��O�F E�H ��c��'`�¶�_�N)�gL���E�����g)�LN9�o�S��0m�"��=���E^��v����'aD��3��p����.��l)��ٶwP{�.��"�L�*Tu�Qu��)�g4%QGBj�$�h��K���qg�r-S���%�+_�/b�������3L��ʎ5����N
� G�yTNWhϻt{x�{�<�}��f9��AKBG�S6�W�=. ��G��7t5�M��Ό�Y�蜵����<E
/%{�x`��̣1Q-N��#wC,Ԇvы�+���*u�m������:["yVA�о�饉)��!�_{���n��� �Kn�K������D�n�ӂB�7ܳV������^��X��-<�j�QK�	-�u��<�u5�U
��!�VYpKf6hD���3`�i�	��JE�%[�#��	��F��a�3�P_�X���%��!�_$Yh����j_k�O<"T��vu`@[eW �3U_yՕ��!�D~��w��D�ޕ�L�&�X_���ެ*�{�m���@�H'���,��E��Sv����t�B�hE�|�t? u^��p)!F��[`\L� (b� zg�f�>f�60��(���߿���I$KZ��%IѲ<�g�Gފj ��D�HŢ.U�9�T�S?����d�D�
�iZ��r%7鎓34�����ʗ%�?�6�`��T�N�b�Z,�{ڛi���G�\������w�vvê�%>ތ��}Һ���)ٙ�(�������*�1f��Ѥ�W�n��y��Bm� 8����5lx�?6�����԰�P�~2�iM������O
�c��Q�|:������Nqr�6C�[�<�����;��* B��w�jR��O�;�\	��
�)�#$כU~��q>��/:c�%��H�_�g7�r��=�
�V?Z|�[� g�tKx:G�Q�K΄�[B2��>#n{Î�����D��@n��jmS�E�ۧ����g1�E@�5E��>��k�u����?Թ�ak.���Z�?2�5p�۽ɆX�ZgBuN �Ap�H ��5�J�iE�l�җ��#� �W���
⥏ງ�)�mL����bn�G�V��P!�R<s�L�j&M��q��Jux9�$b,n�0� �nҮ12�΀{	�B����-3�X�\�z�~|-���];�j+��!��M T��0V�����#��x	�z���/Q��|���]�1%��f�ʚ��=KW��۲�aDT��Iv�#��TQE�-�А�]w��c���\g3ƻΙ^����Bŧ�~h�c�^���:W?}�r�������{�k��f���6Na���Vig?{2�o�0;�ݾ�P\�E�P?.��4�S�|�vaJ=��󁜌`�v��9 2�g��'V�>�-���,��w����{��h�zHQD�rߎ��$�B��������
Y�G�Q%!D+(,���O�E�����
�<Uϔ�H�q �m&�u��Y������U���
[@~}�+	
�G�إFa��F31O����os�O��Ax0��i<jg�%�
W�&?{���WJ�&
�m��>����ի�:��dM�[�̾����_:��JJ�wC���&��	>�x5{kh�}9��kUa�=opr]]/�mx��X�E�B���S�:�R����n�<�`�B���.غ3����o��6u}ܽ��p��9س_�S�'>1lp*r<�J�Y�x)�Wh�@/s�4�6���k1m;��)�����y�!��5�LrV�s!��DK<LK^(�s�e,d���+ӌ@�ת��p�J��Dz�e��WKt5=S�	h�Wc�b��×\��Le�ZȳP��B�q���-�w�g��,�˭b"r�h~]G� �66>0H�g`�<s��W�	x�,�Q�&�*��~��W'�D���:�u^��o)�֨V2U���n�P������=�w���du�3��.�1݈1�yr��n���fr�;�e�;�"��Y?���K�I�(����0!�bg,��h��7�3���s�G�NIN�9k��q�Ξ��۪Я	uD"/*�7n���b�c,Ǚ�,�m�R`G�{]\�ڡz{���<���G��B�����i�׋�|)�_B������s�#W����|��ݗ�Ť*���2V"&Ỳ��J�i�m�eWxz(�&{Y�+�׋�����	V�l�Dǽy+wH7���Gp�1��1<K[L>�d�����l^���fT���{M�W<?��F+��=o�Im^MR�S�G�i4'�莯��#��G%�o�(8$��I�I�:��I�8v(���H�@��<��eĳ��
�J`�)���	O���^2(-�؅@���c��U��T{i�u��_��C�N�G<R4X$ִ|�z�f}:�;���i�$<^hP��\u/^��J��p���1�/��A����s�h�$�s ���I�����a���;�(r�g���巕)��p����Nb8��
�b�˭��h��-���h#��T�Q��,E-j3*��������xՁ�O9��b�7��ǌ����ʣ��R�7n�^�O4�-�$��%��{���O�3��8�ny������c������?�#�Q�kn�x[���w=��12x�JKq~�7$�[��2�9�'ᩥ���d�V@3���Ը��/l2���lwYc��M1�B;���R�c��S���?>���;p'���[�9���C�VV�N��V�r�0	�+!��|���`b���8_rk��p�������{��YL�(`�0��_�ua��������`Z���d\�D_�kn��������D��N������x*e��f��i1�C��[��Q
����_����|w���^�⾠6%�1fGଠ�n�!���);O(����K�=c�C�.�j�*-����maDj��'��g�w�<�*�{���;f;��`��IN=��BYa�+.GTĮ�a���!�-j�L�w�h;�8>&�GHh*_�KD���F}`��C����y<��+�S�����3#����qiTf���Mq�����lEF��L��?>�Zi q��{��k�6�4�b1���3/�4��=����9�GX\4��.:)�X%��{!�\����)��3�A��h%sȜ��%��2�sAC���L+�e�@1*��j���!E`�f��u�)����'�ُ�N�a��[uN���+S�c�ҧ۲��D2.�Aj"H(U@��h.BC)+�c\;dէ�~���L�a�0���Y3l��Vakd{7 � �x�Rθ"h,�r����m{D��O�Y��!#�p��֋�3�"����Is�b&]J�B4��|�'�e���5�|_�d�w�5�0��O���%ܷH�t˹��s��<�?�� e��9���(�YFvQ9�� �H��}بe�͛�@�Q��ϱ�<NU��Ur	� �i�&��:�&$ELCE0d}K��� �]����/��:+3��^s�u�lƷ��f����!m�L;�����<*���E���h=����rH&f�YZX�)���n���^~ϕ�g���yM�N�!��ؽF��`�4�rDP?�3=�X=�{�}��?��}��1�G(�ت#9Y^�;벁�)=^�)�$����Z}P��O��_p���&�6�D�J��}�3�j��FG�㍒��_(��Е�#V�t�r�
)\.q˿�OZ��d��NѮ�E�gL�M0N����CIw�����k{G��l
�a��9�:���ƚ��a���5���6���c��s佛��L�W_ ��"���~���d{ ��)�źD.\��$����#{��1͋�V��� //D�}�2b���E����'U������1����d#/˺���$��߹��4���_R,��J�*�F�P�C8y��[~ �2�5E^c���G��#�|�M�,�9�vK��j\���m1/-���m�$�j��ɣ@ �#�yt�'ͮ��%��~��z��ߠ�I؄n<��#�8һ��Z�&�z��^PÒ�m8���Q��K��z|M&�������=��L�@c7=�{�ˁ:�vDؑ�y�a�h��(ne�'K"����&����d5	��!�/�f/S����t�j-��?�d���H+v�W����V{�L���+�+�#�L����B�^;��>��Yjw���'O�mR�p�x-�a� !`�]j��Ϛ.~���^RnH1��#i!���%Q� ~-���t��!��]FI��#
��+�vDȠrǀF�x�U?���`K�!�)�[���\=�G��N���������&�O#m��m��I]��q�ٙIm��Ϩ�����ǚ���4OTo�)b|q@AMˬ��j\Q����k�$$f^����-1&���f� �����]nu��'�`�!�8hd�/�F��f�_���f	[��S`.�)��j6b�/|����XV]��Wk/�8��p%�^�Y �� ������
A��p+���wQu�$�N<�\{��Bp�68����j�e�֒������>M�4!6�T��:��{EӍ�LB�k'b>(��E,1�}\F�m�ė�Bɿw��z�~�m���	�r.��g�I���W�p��9����J��2�y��yv�dL�;@����>%�	瀟 H,�d�?}������1����1�Ȓ�P����>���M/)c���B뮣��������9�D"芀(0��!�ڭn�ՠ��F�h�.��ў0W��ro��m�����c`�M���#���=\�AE����"�̜�v2z�#^pYȟ`wCH�=�u�T�s����Y]X	j|��Z�'�͘t�`�1���m�D��v}FH9�6��qSv�ְ�-vޑn�-��kVP��c��<���P��I��O��l�U�#,<�:ov� �sQ�����m#q,�P�M����p|�S �z�ȵ�G�<��h˿"@�eΟ�M���'����~s�2Y�h�5kf�����nBW�(�!b�z]����"-�ɤ'�(���,�d6k=�c��T_6ڽ���&��艛�>ۡ��h��&�Y<hAs�oϞ�����ֈ.+�@(P��Gt�ȕr�<k #P��{lV�'�+�qK�)3�[��k?\�Y���py���P�ǳǊDvZ�y�rj��𛠲�&r�Ķ��z�,�X�@w�8��C�.)b���� �B!�L��	��9�R�6]`�Åt^��π���D���+{�\4w-����gK���FՏ�*���z�cf���vZEbן�1ˇ�}��� fD�#|S�B$���Tc�YO�-t�V{γ����I��>���Џ"��2Q��r�ř�Êa�9�����K��׋	�?�:Y��j��@֥]�{�3�X�*j0h������/!b���H$��?X�Z_�EkX�i1�Q(�����l={,|��U�ȟA]����t�C8�Qs����elko[SM`���%}�lTz��������u8S�����I��PO�9�����G�$�d9]��0�����c��y��{���a�tL��r���� �8�f��~�u!`��8B>V��.j���"�?V�r�[|Ӻp�J.XK^ת�d��.�l(�6����k���u��v��^��u��pnm4N�R��9��+�0D�M�Ur8��6�,	���)귳��8ʅ��8�V�Dҩ�������R�J�"Tj�]��a~�[!��z��"�nbg�a�����dx3��u�����b	TG�28,+�|M�������֪h���ܿա�*$>��=�O%�QcF�U.o�ׁ �s��	_N�����|(�6�Ew�������\Gu�`Y?K���2	V`�\�Iv��Lq�ZK8b9E�c6�,^:?���Δ�����6%9��6*��\��r���zs�SE_�v,���55���UD�N��(���^W���ޜ)�֑`�X���v}N1]�g��r��I߬��+?'i��z��JV� G�L��jb��nG��v��㛽]ׯ`�@�in$�[V�W)��f	�Z�l���lII�~��y�Q�T_�oY�.6S-���+~Kq�]� 4K�wQ� ��޼���q���`��".]D=3�,���������|'��+��<Q�Q�ӻ�W��SrL��O���<���
s��˓�GƮ���#���H��O�t.O���ɧhKP�jm������0�7'�z�[������l�۠)*�b������ٷ���P�`7%y2�Fխ���<�ܧ����_���ޘr��o�"����Ȗ��\�u�ic�'�NB��N�4�)V�~�}�Ajcd�b��͠u1�ܶO�I��L,i4��5K��6l������\�P�*�2i�@rE;��:���cw����R;��1M�'_�!�r0�Ca��h��К�j��E����_�
��Uǡ���V��J'Wv�^�ud�>@�� я�.](sm�n~��EJ� �W��T3�-�M�n��ג���U�P�VE��$������6�d���,�H9�V"醚p,+���l�T��nD���,(n"�h����Â
\kU���	1�2C��0�fg�E��Ŵ�2�ح�G�u׎�gz���3	�:��P^� ���"�h�"�F�ި诌���wA)��A�s���2��7�,�>�V�wr��J�v�9#ϯ��L:���/I�ֽ�=:�G>�Hgr��������S�k-�� �U���8C=@�f�NG��zԠ�DE��ߥ���A��{���S�a�5��n�l'�#	�3���%��~R��I�,�9<x�6�0Y�8�\��A�#`�����%P�yQ�'⼡��t�� W�/��\�L��u�Sf���V-�r~�2�/��;�%���-w���Na�����'��_�g*]՚ v�\&#Ѭ�ꑓ]9������q/���+�ů5o�� �=�n#��R�^�i/�#�d�y��@�Q�eЖͺ�pº�,O�z���&A��{�.��]�^��q�$��t�b,:�TM�y�b9���>�m	�������>������i`޴��8j��e��@*Jh>����t6
���>�LZO���a'�{���%Њ�b���zf�(׉�B��ǂ��mB���^��,�Va[�����B�_�쬙���C@d��Mg��P�N4;���:��-'�(�z�{ƨX�����JAZ)�4�o�D����}��)�Z�J����5���ɚ�0�u&0b��)a�\B��vY�����,3����5U��P��H�U���/��o5�+)������]�|���>@h%�\��d���8�Ll��;��FV�4�@�W�e�e��
����g$ak:�~�$�����j	f(�6*����z gM�����'g�U�(D���?4w��8�P����w�$���	�(��< �wa0<�b)��y��Zq��`W���f�@0D7�X���7����Q���T^`+�Ѐ{J�`>u�N� �,��y#�>U����Qh�I�J�)�l������5��VA�t8�����ұ�2�g|�.�@;8Q�Ж�ox�ju�����U��0Ʃl%�v,z���Ѭ�?	s<��w��9s>�y���L�c�V�d?;2����T# "�g�dB�0)$�d�\b�a�s�E5K �r���8\��C/����Q���7�Q��ι�;�����'���Y�B6t��[~2�p�=���� 0���+_nkg��ow�p��ss��B��^|�j����ff��@(>�W�4Sq����j���.��ת(��&ۄ/�M -�~A�cmԳ�/�~���nfC��2�"A> y���`��?�P�S&y�4_;u���*;�ق]��c��(t����*�(��x=vz�v�S���qRk�4vM�jkZ�l�<3G+����>m���#eӛ�X_B�5����;iO�֎���u-���)v5������2y�4�k�28mQ��6���px���N��}Z��#��O��ί��4�.�E�L���,ٗ5E��xQnʕ'TD~.����yA��yġq��P�\�r�/�VXw�!��¬v����`����`���e* t9�juIk�t����10C�ڶ����!��:bK�Q��o>!7�Tr�)|?$xU��'IN�6�Z�@:^�{�J��{���-�}Q�o�}r��HL|<����*����?������b�����t���"�:I��+�SCCR"�B�%Q�-�U��t���/��]d؂�,wт���}\���@G�j�L�B} ��,o�?��M��>&�G\/�1qk't���7P���}~8tf'�r�"f&�O�7�X�Ӕ�ϋ�z�r�_�p^�=���S�,�&ңk,�55������[F� �N5�%��4�h���, r ���5��|CJ[[z&�ؿt���*G+�����|۴�~#�T"�����'q��1��Q�J[r�<�&G�����Y�7������o^O�p���^�M�R��a���do��������b�z6y�h�=h<�Y��<Y	~tr��U���@�5�
V6-wS���(k:xLYb��"��K��1 W�����=:²�'ڀ�N��.l�E�w㥃 ^�X���w�0��*H�)�| �����0?'E��/u�eS&p�*�� �1�x�ķ}�eGf����س���j�L�N� y9�"/�|��-j���G�yi�e�&�e�i��#�P0��$�^Z�N0ݨ$$96,�@άʗ*��O�Ec$~����r�$هQ�mB졖��hE�����{g[wT�@�Bѻ�g� �:����N���Jv�kYb�!�eb��.���4�����vr,�,�A3�*ᦲtK4V�z~`.����!�t�y���`�1	
��$�&ׁm�T>qb�������2 ������8����4�|�oȵ��[e�JI���R1�<��w�#�6�vd:��ŏ_�=UzM�L��dhyyU��H�*�io(To�f[�*9��L. �X�E���u0Q���"�N �Hwؙ�\���J����4�j�%J�S n>����Dx.�P �J����+j_>���Z��9��~�!��j��[�'&����� (<�-�
:�F��\���w�8Rr jr*.+������~Y��$@�/l^�9�G�JRo��ָP�X����0��n�� �
�ݢ�����GD�@�ur+��1�i�Y�h"��#�+�Y@!+f�9�`���ޒ�I�~�?��¸��/�ȕ��}i������s
�OT� �C_��.J���~��Α�$"���#�����?�=(�|�Y1F�|� q�%t^����W�n��Ç������ Fam��aT)GQ�x+�<E7YO:����z9g�ůsd�8��r��v�,��g���"A����j:�k�@s"��@N �(T��r�0�4�IP�k`���r�V��<#��_TF�az��<cX���N�	��|;�ZY�fF9).�~t��H�݁�8<M���7���C\���2"tOO f;u�s~]D�?9�bz�*\�O�B5���u�L�+(��)���cW��*V�U+��Ӟ�}��)�߯0�r��-Xb��ni@+�,랆-��s� a��4G+��^�j��{,��-�XL��1D�;v��� 0Ԕ�$��+��#r1��Iѷ�1O)ݐ@��b�r1�x��� �}��eN��X=�j���n`�k�}b)dÊ�d���<�=H�!y��s��s���&t[&1E͈��v䥡�V1H�wwW��q�7��:��/��Y���\��;в�eH�|��k!�������d�-���&ƾ��n���]0d�� ."׼�d�wU"���Ǡ��3ũD�S��Y�<݀�5ŅW7Z�}2�d���G�����ސ����xs���A����o'nʹ�cGz�o�8R:U{��z�י�����"�]�4�etL��qC�*;-�h�ż�U��Wx�U��0����R�r��}�	B�p!��5/2T-�1�_�j� ظ8"���ܒ�W)3,u�B�"j�C�p
���-9�hZ+����i�[�`�N����o��nVjIg�кG.��"Foڋ��ǵv�>œm��t�M�rNi�]h���,�?椐�n~�k�(����W���ưP���s�$���y��u��N<a���B��aK�^�r�T�A*�Q%2[���<�?����C��\�Z�ї���&:c2��zbxp(d��X~�N�q��$kw�J��%8vٌ H�3��Y �:UA� R�\V�*r�z��nB�h!��-���j�S�'�D����*�e'׹��ޔ�%�cs������B+����p�@��R�?�ѯ����ZU�m�g��>Sr���������h��;/{;iD� Y�>��)VI�w��}�#��gO�Iox����D�R�tgr���8�'oZ�"�T�Ll�/l����a,4����m��$���fK-b�nL����v
B�dt�>�u�8C
(����Ǩ�����Ɂ���n��o$��]B䦐�?��!,���DC'�`lO(hG^6c��w���V�����xLtoS(��ՈOAA �*={Ō���- ��^���9��FBa ����~����&���[YAb���1lC|H���In�֛�n�Z��˵�<�6>Ȱ�Y���%�2USb����ť��K�8���ģ�X��|q��f-�N�Z�w���_"q��Vhm�>�*��z�+��P�^eD_ڡ�v�e
q%�d��	R�,�����=p9��ܼ	�L�:��Dz_d�JT�6s�
6�+V�[�<w2S,�5�S��bY��/LH�5(�W!S$ٶ4���@�_�	Ai?I7�ޱ{��=�>U�.�a&��|WO� �]�'El������l�n9�8t���W���+��&����G5-�\^���3UA#9�̬��e��i�\TM�iHg���	�y��S#o$��E��5Glx6��	m��ߐ��J��J��,�>?`1!N�I����w�͋ ���*��@.�t��0�^{�9x۝��Ӭ��X��@!ѤL�b2׻���-�2)��QF��*�:	�㺊[�"B�g��L�<�k���`��u���f�x�]G�Q4��4��C>�^��Ղ#�{jI@�C����g�!�%ޮK���ֻ�ճ!&�g�N��Xp����qUU!u>D�
:A�9��CXo]�g�r㑻��Fv�h���c�}s�_
��g�v���-�P���.�d�;��d�4�nT�3��3�öf�N�țBc�Ȗ�3���g�-'�g":U�Ye]&��yxӶ�&&B��e��ɟ@���I��&�GV,��3�z9�?@�
т.D*�*�F)�������
�X쩠�{1���X���;@9	�&��܊}���g���q��l]�v�E�Ht��H5�ďIb����E6/�mV����L��B�Z����5z�q��k����/�ڣo���),aמU����������g���1�����g~��/,��j*�E8���IxcIe�E��LR~{!<=
��&co�_&Qk�[0pݫ-9"xד�L�9q�1�%�h�l%9$��E�h��/�x�}����zH��V��_6��+f˼�X��^F�N�3s���_d��������w	������4t�ʖ�P䟚��v���w��U��ֲ�{O��m�7@������4p�5��aK^���
B���0og8L�V�q/�.~�����a+�嫖AUPx|��sR�C��8!]�W�]d`$y�cޥ-��d���-��X���2��h4O�3��J
���������θ�t�U�y5@��s��@��g�%���%�!$�8U��o�Z�$S20v��Fa'��d��D��փ��E��G�5�/�/��=��v=��P����wk��ٞm� [�S��l#tr�e��~�(��X7��yZ�6�XR��D�ǎ�V�� �
u��F�z��0F��(ٯ�Aaf9�r�ǳP]��x�ܽ������Kh*��t�����DFg��3��y��T�l���
!-_rE�*�P�ro;�J]���_D��R��JZ�U"�0(�,3�2��!!�0�Z�~k!�9S}bQ�Jp�0k����bQ�P���y-�}.³�z�A��BV�R��U[��M���9G������`�1-j�s���a��W��pX�y��i����@?��jK��j�����)�C��_7hχv�ag�t'��U������+����͕Gߴ�LW a�3��[�A�@�"�|1�rb�t��N�>{��z!��@����a�4�=�6;��
�Z�x������y��YL�y��#`EJ���'�4sC�U��h�4W�[:	9 �A^J���,����ٿ.��ݕ�����5�j\��ͭ�r���@&��9�U�4I	i�J�M@�H�P�G��b`�i������# )u���Y���m�8�5�m�� ��jβ֭���_�lآ�̓��Xi9jɡ�B�,�#��W��]U�~�R␠�ʥ?��}����ZI� :��dHɔ4�����i�xY��^������Rs'�{'Ҵ���gE%1��<,}�Q K�w�⍣ �8q�8����ۊ=�;��F	KL~/]�9�G��&�S�)��~yN��՜`�6Rψ����v�@����������>y�:%LI�.�{��Ⱦ��la����s0Z0j!^9��-�3�F9�������h͌Cj\��Z�;��v�5��Ar�Z�$��2�,��
���j����t3�~(�^;�c<�.e�Z��x�E�}P1;����L��䒙i�{�#���D�I����ɘXʡ�Z�5�C�Q!��W�	�a�)��(��E3EW+k��)H�j�,-hk¬��4$d���{`n	F�7~��DC�����6���f��҃I�q��8�l�)+"ܬ?v�Ծy+��U�����H���~^ܚK�li���D����2Q}�E�/�g�W?���4�"��OP�D�۴H^�ut����s�W�Qʪ�ʓJ��*��V��"�2ڴ)N��knAu�0�ټH�,�q�}!����'&�V���zlSڈ0#� @��/��R���X2lr{`��SS�0B%֙E�R��Å/{q�ʤ~���6y��	���3�M�j��;��IJ���HS�e�mk���+�/)����-U��\43�2"}ȳ�d"��} ����F+J�h�'I&D���Y�����$W���6�>�	���WZ����r"�!��������1����{h��'�u��o����ۛ�JͶ��'�r��wl���=��s��qf��g�2�d|(�y���tX��L���[WH�]<Ot�b����(��?0�SS�g(cQ�a����Nds�|��T3��b�����>UBD@Ѧ0JD~�G/ERK󧨦��"�;��6�
�<p޼����!H9����\fl���={��԰"����
W\�l�K\ {r7�"(�A<��[�9N�5c�����E��Hm	/TC�r�aJ�l�)�5�;�U�CSg���6����x���t��
�� ��l��b[M�3'�@8�#<��E�p�B�U��	M�^�P�(L������ָ|fG�^���d�!v�9�wI΅s]�gvu�Zl�_�bq���0{q]��؄�,T����yT���\�Cq �O�(��X�Et[��k\�#���P���Ur��rEx{��T�r�d�C1��Y!j]!l`aﴧ�'~�7@�3�Ug�5Ɂ��	�MY�P�S�����ҥ���nc���&K*Nn���X|̊�s}+���,�����,i�=����(�B�)KT�J2�H���K�|�����,��A�D���:�|'6y'"��Jl���1��0����E�X�C�f6�]{L(����OΆ^R9�����=��.q���vB6�Al�#�ʟ��otD{��uٻ�³�0J��|��K��1	 $�+��۞��Ð/r4�C];k�ӎB�olK7֞!~ ����s'D���uuTe8�A�8/��a䊃��f�7v�c|�N>K2$�I�/u�>1�!A�C�����g7����fk���ȞB����9���ԬX����/S�}����fѣW�f�~yd�t?�X,�x.x�̗H�d)I�
����"�ˏ��2��������u�����8*�Pc�j1'�2Jt�˻]S�Ny��"����qo���g36�$Y�p��nOzT�F���D
W���PK�Zw��v�t	3r�d����ݖ�>��[ �&uC�O>�k3��������Îun���7�8q!Ix�h�Y�N?�R�8N5~j����3KP�2��tr(�RVn�ꜹv,�<�zB�ӣLڝ�A1[��vB�5��H�V�q�|��� w{Bk�8~1.�Hy��r��&D�ṳj�|���^�D��b2�s��#)����k�Uq~lFYza�����s,�Ծ�⎈=[�\H���y�!�e�G,��i��yвI{��1l�H�kvE	r�.�*�oF$��Q�=�J�JjfO*�n����Ε=q=�(�ߴ`��8�y	�珆�'�B���x�:j��!�?T=-.�X*8Wq���X��)�;��*�&�L����b��o��Z�n�̄�4|$�zVv��
9E��aP(N�4��W�*�v�'K$�4�:^���ߎep�f?�=V�
7u����(���(2Xe�o��c|�YHR���������<�_5�/o4g�&�����f���C�����49�/�3�Cs.�:�*����p�R�S�!Ϣ�݃}��xc4I�u}���ݨ��N�كDJc����t0�_�r:7#G���C&�.�\�Kh���r��x	�L��Yp|�� DC8Rs|�xτt�Eؒ�8��D��U0�W^7�걓���8Y���O��M2��vF.}%�އ'ࢅ�N�X舗�+w�&IVh�CϚ�}Jټ�-dު)�pE2w~;.���.�U��mPYnL��:�G��}S-�#C0���=ʷ69�e3����H���:T�� ��4��u�ѳ -T�7ȀW����qgp�q�O�_�4]7����2�÷��*|C�*�B�BU�˦�
�0�_'�$D|�2݃`pv;�l/)�r2�+?U\��`�X�r����µH2QSc\�'�Tբx�4uT�wb�}L"�$s�|��E�8�	�%π�-��"���z7�����=8��i�i�Yt$,��>t�DûQ"�]�Z�B�mn4�����Z0��\ӔK\\�f�\Sߞ���D�c�4�����H#���"�>����\8�o�D���4S'�^�'S�b�,4���y�wG��g��	��Ъ10��7����=��V��8T`�(\d���	I���E̳H����E�g��ɑ�6�yOꁯ�\1��W1�֐S��m�R�h-�>i�����Ys�gZ!T���Ί����I �4�.Y�SR��|��LoM�)XG�"lfh�j�Bg��o$ ^e�r&"f�&������M�aS١>�O�M�C�d��@�;%nhy�y��IUVc�$c�i�y�j�E}��P����WN����P,��U�D�)w�g���N�>�	ވ�x��p�w�g��r>�0�E���@�Ft���j8ր[���؜ j��9���$� �R*��#�N}������D4UnB��q�tz@�ۀ��-���KG��I
�[�xT���}[��g��x3o���
N-%v��U����%�5�*�+u�d�EUH^�\�Yg��Z�6z����e��_�ζ�ve\��i��>�cg8�o@�!)X�����$��I�q»j�]Zp#r8(h�O�yS^��Ku�����, �@��O�:B��ņ��"�6o��t?��uBL�eH��>����-��b�4�pm+Py����ᳮO���lu;FÒf��Z�ֽ89��-'��Q
Y�`��g;BAk�;	I~��}���?�����"=�'�?}�>�f!e�S�v��*�m���en1w����K��UMe��:p�q���/�3��J~��RU/yS�i������1xe���l�W('��r�(�%���ky,�d�J2+2E$,&	
�[���>�_Ŗ�L��BO)e�&/�	�k|Q<*�+5?VIߤ�29 Ul�?v\u��|��b���픗�N���!n����E:G@��a�, �;8��Isn�5�9SʍȬT�z�cQi��}:kueS��%C��E{�� ��缯�+?E�u�+.�L�:�K��L�1pP�Vd���/��_A�� AC�nYOK=������0Q���{5��87���zI�_�eV��F��t�op|*�譖=^_
�S9��Ǡs���
if�{*�����?����[��u{;EaX(J�}�Xv8���֍�/@���JǶ�sIs��Z�J�����d�_��I3ȃ��,��	Ƹ�nϒ �P��2���qc��d�o�PG��'\@�m7{fF���T���!�6Mq��]	T��/�w9Ԥ���[c&kXM��k��s�q� ���4{�����`���<�FM�CkH�y����!����6���A2���]HSXB@|��'��D^
mo��YG'2*/���Й�������cz,���5�І�:�=��VG�\�
2|�W&s>���	 �M��?�)������H���<���xX�7B�t�9A����3�#v�$Y����	�V�|�^�19���h���i�(�
m���f���s0!�RT^fQ�m�v��wX�&7&Z	���n�\�
�&�P�?n��jCQ�f��b�.gAy���w�z�#-{�`J4���jqv�EN��O}�m������)Ry��B*�?�z]a*��((�墤q�`��S�A����od���oRŮ��&ʷ�˻�d�KzFAb���W�q�9z|r���+A�y��Cч����ֳ��F�Cޓ���>0��*���6��#�\�(~�TGrm�V�AqyV�y�EFro���qBȗ;)r�*f���S:Ӎ�i	H�<M*m��s�.�CN�RqY`S��C�D�b���o7�Q�;��$g^ ����=�Ov�|'J-��M�C���T�nR)68���PY����Z�#9�B�9V�F:$2c�?jt̿���Ǒ�с��1��}o�6��'�C}#��W�`S�������1j�0f|�������p"(�讜�a�5��֌�X�V�}�b�N� ^#������m��66�/�]�
,6�a�_4�tu��b�3��*��hZ?<��1�~q�'KyS��ɫ�1��E��)]���,`�fn��V�$5������b<}�t�6������Z0&���!lƂ�vӚ�g~�����5��B.�z�A�"23&8�ʴL�^�)�O�ݵ=?I�����C�9!f�a&�%�z� �/�^��NZ��;�t�G���A�0E�=ةD��|2� �Q��ӣ��e{�v*z�B��$�~�<!��O�Ju�|J+7̩Q��������m�\/2����ŉ������)��e��?�U�'/��$�5�GȲ�:���ؗ��P�^�_?�K �oAR&l��R��<�w�����ZK�m��*)�ԍ�.�@��+/�sq� �0�uS���R�	�i�O��o�$w���,(����y�[� �[��̰�ZX�\<.m��!�PÑV��)���+����Y�##��H{�>��Zv������6�������"�B�xB^^t��<0�7��aOά����2������`,�����}��������|�g�Ֆ�s#[.Y|zG�NhД��xV���H�Z�Q^��%#����� �Rl���) �G�J�)A�&�H����vS��."�mrQ�';��gH���} E�Oh3��ݘ�ju��Wg�a�y/A��c�8���.�L?j[�*ys�=��} �#Y���(m������b$$Y�h���?u���V�g&�h����\s��#"�F`��r�D�CC��˰�����C �2NWq�T(�&x����(�S7.�Ɖ"H��kE8=0>����#8���'n��ȌP�C�F�,��	iCy]�l�09���ڨ��q�Ǫ�b����%u�*7��}�V�oo&�:s�)����s�� f���f�׽�mդa&W���))�6��Y�,9��:��!%����HHbw>2�S�E.���B˸����C���bz7���s��C�/�&�M�a�����Y4������P���@+:V�Q���p1.uz�ȤX�1�Z����NG[u���{��^�du�O?��d;�`��vpb.�4:���WC*͓���'&� ���d��	2p���h���{G-G�W/�$��֌I.��ۿ6Δ�̿w	>~�tУ(���1�J'�M\[��p�B�t>}�S�������+�Z⏊)V���k�;�v��md.��İ}�d�XC�6�T`�Tw�3�K>��b�W��۾X"k�`�Xo|�f�b>��q����-�P�(���S�p�N�E���t�"�|$`��څ�I�T���Ԑ%ú��5�*TE����-��"ޭ;���Y�6�
h� J�ӥ�1|blIw�`qn�R��O�tD������EZR�2�h��	jP_`��*�0��y�|K����TFNB�n�=��V�G��	=��>\����:<�����wS�<�
���~�ه������y�$�)V���$��f��A�X�Hx��7M�o?-�T���
r%ѓ���5:�_���#J|���F��C�ͯ|� 슊�X��X�RǼKy�3�Qʀ����z"@�:
�E#�cz�*�
Uuw!h"AA�����Z|�
OR�yx��R�K&&o���2=x)��+��QG|�Q�'���;�&T�O5�J$��^���4Z~Ƅ$֣�:�9���M ���s�k�bc�2�G���c�����o�.���f���o@�8Y*�����M��_gD���x�WBM��m9y�!�^� ���9����Hzo�XK1 y-TSV1�jս�?7E�Z��u��Ԅ��Jg�jhP��.�$�TY�FN�8a�ǂS���Ԛ��y�(�ab����B�'2�
5�@a��Ԏ��`bQ�j1�{��(��zK�/�����+��o�z�A�c񰘐��Ǖv�D�ڤ�aU�Ӳ9X��hgﲀ�\z ��b�ݺ��gŽ�B�����Ͱ���h�S�yL:�T�,����?��$�aG84����o	�~�/��o��'&"�����%<R�
�{XI۳Piz!�erP��$8Fݯ�L��P�����W3��#I��µQl�;��mz�21��8�4>S�2N���iS��a*��d���/��!��#ΉN�:�>;����m�@��(+����=�(�(#ړ̏��۪(F�zA`���AüԔ���������I�;���-�E���\(=����*�P��_�mV������@�?�Q�4%��.�d��b���m�Psi%K֏��.e�A�`4�&ck`�x����ٮ����+8��@��qF�Y�4����Zt�[F�����A�!�ɴ�?�;�#z�1�ٙ��J��
���	Xx�?zN�Z.=��Cv�"]:�knP����^�d��˪�O��ӓn�'�C�/�N���&�*Mf��IXe�ms��x*�������Q��Z=W��k���ŶK{+t*���w찕q#6��˔ /M��0�.6`;XN�E ��9;d��
���p�2I�,G�@SFm����Η0{ rպs�����j������y�E���� �_���v��~PS�i�0's'��ʻB�����4JWE0>m6� N~�[`>蔑Ӵ�ZM���lp��2���8�ϲ�ū`����Cۢ�#�}zO��H���7����b"2!ѫ|�6=[�Z�m?r�$���/ٕ-��`]�$R֢vf�<E�}W	.�̕�+�f�a%;x�����>b�
�F93T�G�{`��������s��?���=��)��5%�? ���Bʃ���J��ŉ}�w:!�/���\���؀�ፓ[ڟs�F
n{:ߊ���_�I4��/�C�)��ڬ)�������g�0�wܰ�Y���đ��:Mj'9�M9��G �\1ŭ�I�S�;H�@R#J9��g[�~)�oρv�b�O�����}���Va�z���>������u,�.1�,h*���VӇ��훔�Net�o�@���M���� 
��/.�BY~I^�j��S�����'���#a�}�I�e�zk>:��A:{���>�b8�A�G���8K�R���i��K�8�vn�c���j�g�S6G&�+C\�b��Co"�ήU�6Ώ[�`�w��z�0����R��I��F~)>4@�]�#6�$;t�u�Qlj��+30���
kp��3"@Nm��i��AE)��~���snKU��<�����S�qY#M������՚Q�m�!($Hme��b���Լ������o�b�Ag�y�jBZ��F�*\�Kd���uR?�d�J3K�Slºՙ���;/�KiZ-<�s��L�%���T���m@�]`�\����LA�꣓����ˍT�(����YYf�>������?��r#ԁ:�܆������,�(c��_+��
��7?s��R�/�Y�5�$M� ��0�	1c��q!\��/0aϞ\�U�1!�c�T�Wz���?�3+=*��Pw<��) �~�\�����p��z�gmӷg�Tc�j���:�2r��� �8���4n^J��C����d+zuI@s�+�sV(�c�I7^4��`�B�Y4��Șo�&0�J7}��|-��^�|\5)�����3�->=UfB�|��-5w����AC�k��u\�#ns�jz�2���j�Zv5�7@`���8�ʼ�|���`�X��I�>4-���o؀�oj:*�]�]������g���PE���"�,�%ap
r��Q��A�H���T��A��K�r�Ug��}ς�'�RŒ~� N��`ˇ|�QY8���A5�����U@�5�X��)D�-'l�x��&���J�ʥ��.��JH�D�2D�? ��ܦ�И8�L�C���調#es%��ۅj7�{.��p������G��ݏ��]v#��B�
��@�C�#}`w �=��,���K�aY�������"r�|!gd�%2¾�wˀ��d�F�tz
�ѐK��z���{���L?pſ$�@Q�#M��0u���m	��0r3B}�p�|v}�����;�����,���>P�5���U�שc��b���NWwYA�ύ�+�S�Vʥ��G�R�V���E���O�1��Y�o��=�c�m��h��5��g�¶�F43e�k���=�!�
;{�1%!�N�~yo��)�p:�<��"�:~� 
�#*�u@/�I�t_���x�r!��R�GnZ�I<����:���H)��6rd{oAg�@ 4�,��%���#�W]�A:�Ew��&�uҊ� �z��Nts�/�O�5!�)N�e��W.���J�:9̒�8G���\g���;^���=q�|f��ٔ F������T �I�П:�N9�Ξ��cSape�1�.a��h5�z�<��Vj�7����Ƚ3�
o�x-co�o���-|.P�^����i[z���ZE�!Ҍ5+���o8�a�N4�vD�t��_��ȍ��Һ�3�uL�W�c�ID;ySf�8�0I��X��／[r��^$APΜP�2T4�j��t��ڥ)��`��d��D�D���](�y=� �BW��ج!؁�$i9��)r���UP�?ī���}�r�Nk�YHz�\�m�'<-S6�Z�w�qi���?M>i���H� �����pR5��<N�òn}�Ă�A�
2W���Yd�U{X��WYXдgOή�0��/l*O��Ķ������cX��ŹL����ll�"�c���{G^^� �XwV��?p[�6ۂ�7�Gj��Z9vRk)ԗ��k(((�F7�Z�BB|��[���L]��
c�L�����q#B�
΂F|�]EI��E�M5�>]ֱ�V0?�	�ZJ!.���P���tϻ�G�b��w�=n⽖�'JLm�F�#��{��Sp)��r'��+Q�~jp�pnqs{f�P�`��p����c;�z���� �!�h�i`B���qZv\)%���V3�B�/� �`t
��?���^�����ϸ��.D^6�Qiw#��I����\�v��T�HG5�F����U���s�"H(��H�Q�OA*����}�P�b�6�Ų���#�9��ӚΑ@u�1���\�
�
���1@�t"�驍���N�$'�| &J6GF�|��j�,n$Bz�eJ�#ӈV�v�E(�ǒ�6t[��#Z�^�� �t��}�Wx?F��w�|Tm2���*Ih)�r�2��s� ���|�� a57~\Ǵ~��^�_��v�,eY�ˉSh�;P�&j�C�,����}� U�y�9>03���:�S1�k&a\�����]���	����>a���'>�3���=���yL����wہ#�D)�Q�h�ߊ� �BYU�P�ᯄ.-�˟��"BC=3�綧( vNP8	���P����I4f͍m��%�{�I�Ǘ�?o=���)�z3剺�����!��O;��Rk��7���X��S˃���R���a��?Lo\��1� ��5kP;�A���E:H]F���S�M�گC��8~l�|��g*��\��O��mrJ2�ݏo�N,���0���;2G��t�C �jH�릗s�,0����X�1럹:3q1#�U�kl�"?�G�5�T^N���g����csx��e,�c7>��H�bZ�W�6��:/�b���2���Y�����~��\�Ŵ�EQ�pMT�\~�[�n���ס��^|�>�����3��9%Ѡ�}� ��8�B��P�'e�@�u�ś���jaH�`N�0h,���m?�~9��=X���NzKj<�NP�Z�E}!2��z"����
^2e|�XJ�G"�w�ŭ�
��$��Q�W'�M�6�)P4/}xR%�����0#UCK#��!��E��.���o�	��������q�D��IѢ8Lb�i�ߊ*Eӊ��Be^?��@J$UfTH!w�'b��Ch�U�6b^0��%n�b��Df��~�U)�g��'ce�@6�c��<��;�v/���� ������x3(���	��T�&��g],k��Bx�gr���+Y���k�կ���(*r=� �2�����Q�?��[T2q�'y�R��S��R�)�-� 5�~Gb� R������@pfp���M��X<w�/�^�sR���±#��c���C7��?R'��|�z���x;PT���E�h0��5��y�;��fn'�������Ax�+WNK���b,>��,��#��\s�9�-�-���XK#�� 
/���Es�u��J�acK���7�OH1�����\av�vq���F���A�c����j3H����Z�o��'W� {���u3�X�g	���7�PtV�ICd�_+��:1
c�qZJ6��l��9K�k�kF~XV�ç�\�J���rֵ\!�3����2��
��eK�
EL>����p�d�r�m���JA�wX�UW^{��(X�AW�@n�+��H?�3�&��Ak�|�SH�����&E��,L�#�5H��k�b��,��� zp;�*♙~���#b��u��# u��rK�YĠ�yRD��;��#��md�A��*�_���H6'��<���7�w;w+}�;� �E��.�&�*߰��[�۽bU@�����aN"�pv����p��9�nf�wEim��8G`�MH��o�p:����J}�����������ë�~Z�쮝*�����k�����g/N�v�!Q�/���k���^nR�R��?(��а�.cem�6cL��K�.�\:#5����P�O�(�U9�kQ���%*1�J�?أ�G���%��69��v����!�L���.[pE34��I����>��?7��0U�#Y񩫋���ݛУ���@��;��޳� ?��T��*R&Dlm�]�x�i�&d�a� �.o�W���ӥ���T:]�Do���N*Y[1;�߳X��湒ȉ�*���x��7HQ��4J�) q ~�CM�����p8^Sh좏���F��~=p����Z"������jI>�*�A�D[HdԂU(�{����[�:�(��ق�!���bѓє�}�(RDT~낒ٌ�>�k}�Z4���֜�ԭ�I���ss�g������t�쟊�4RP��Y��Ky@Y���#�qF�#���/��I�譛�����u���zJ��ѷP��O�?m��ؒ��5�8��z�*]Z���e�w�;UOv)��%`&&�Su����8��.�9���*��V}��]�m����&�Q�7���0|��L�����Z�'��z&y��
�>��{����u�A��d?�� o�wXc���H�ps�b���iD��u�Vٶ�Ӥ���$���������3�g��|�tF˺�0�ڗ�͝��:��y!E0�R��OZ[�b�Y �%[o����?i����[�2A����;���ٕ*�=��2f;���0���ߖ)h;�5��`se����6�)��Ξ6�ʍՖ`����
�-��|k8��8�8g�۞��!m
�*��ބ]��Q��@IVD�2��k�e鉏� gQ�� �o���F+[7qA(t�;�.s�ۥ�$g��g��ո�E�<PfN�l��)H�}E�^��{l�����u���%l�Yʲ�O�����l� ��f5P����2� �|Y:��Ȕ��h?����o�e���}��'� �rm`u�m���T| D���j���m�c*�7V�ZH�xS�g��4�:�&Y�e��md�#�������y<g����V����Q��ڈ@z��ldV�*g�+�N6�t&��?`�%�ZJ54��R�Af��O�s��xT�jK�y�`K�� ���	8�{5$ݳGY���������K� �S�]�ڌ�%9l���� ��ko���|�lt����#/����W䭝��~д]J��&=���B�CKv�h
���eDʶ��(P�����2wkb��\oj<G�%h������
S�if��� �7�g��7�i�y+[0�d�����w�]V��mC�[�Pdf��}*�X����1�Y��w��mgܦ����e�̛�帉y���4�c�5w_��dq�0���-.M��K�P~G�C��)G��o�$�M�w29 ,_�4�WV�u �X1�y���sn�c1`�Z1!���-`���'�z�Z�"��A����=�W+�� � �"�w�0y޶~>S�6h�0t=����?C��塐�12�2���SGIHa�z����GH�s��ܟ����! F:Ƕ��d��e'��|�����K=L���̤�T-�����z=��Qij�ߙۆ5�h�S������ ��ʊX(#�+��?g�;"1t �Vڐ+?���{��&��^q�F�_��a<�Om�(D�����_�>�bĩʟ�ov=я�-���4��qLp-w�#�6�E����`k�1�asU(�)Fͬ�L�/��x2t/�Y"�vK�_j��_'��7)i�v�&��7eޠ���F� ���ͅ�X�Z�@;��N��I�y�;z�ƚ\⬂��q��j��e�j�Ϟ�R�*A�'̆��	N&��ʎL�1�&p������ԡT`��w���k���y
;��3$2�A6���:g0?ZÊ�
]���]��0����=$H���� ���P� �皴��n?�L�����\b�p	l"��&(clze\�Nb�O��g_��"D2�.�0��/z�(�ㇹ*=�O?��~�mz�"1+Tj��
��Bc�q��`��2�O�qA�іn�I�]^+�]�K'�'Gǈ?m�j8��Y���%���g��q��K����K�3�O�1�z�0�G�
 5���A�9	�U�R+�����W�& ��aӦG�^�6�EL ��`�@ܵ��L��8��IWbﱸ�D|�Y��+��aw{��|s5<8euT�&d�b6�DL�^앞�Ю�����#�r=e�����f��{�n�����7��&�9���:��ykR����5o������,E�(���J��=9H������NT�} ydCƩ�ߴ-�f"DڌB�r�J��P�+��#��48ƮI8��^�G�^�3��K�ظ䄿�?z�_H�e�%�ô��M�.���7������ȩ�ܖ�I`�q�=�c̲@R��wpP)�o̻�����ei�Kt�,�g`���ϝ�>U�Rw�������im^%hDb+�������t���#B1g�k���GЃh���q��~H]1uˋ2�T�粹hD�wą�$��8��ɗ)K�|�S�6��s^���}����zA�7Ifc�cC~􈉜��� ��Y&=d���x�4y�4�6PNW�do�=�x8�e�h�0j���5+�L.��z��S5�h��H��6>��Z	
����x���[$�'%�T(xL<�V8z4�!aQ5z�r��6N���=I���x���u�Y�̪�����?"�]��Ť�W��$Ct�^��`֎��ȵ����~���n&� }��׈�N���,��;�d�2#�)ګ�y��|   �?���e�Qҟ��nj�Ե�2g�4�!'�+���_=��oe�~XL�06��16��쿵�p���+^4�_�����Z�J�'����?ζU[��!�����{�Xg�O����f+�`-��m��魉u��}P�?5�ת�"�`$�������I���*O��м�oo�xr�L���J?�Q�O��qW.F�z�\��T����_ܦ�W��@�H����3E�)1��ҁ�%-����t������R�"fa�y��_�T����MG8����I�(�@Q	��p~Nљ�\��	����i⭫���O�ܢ�$�k�mR�,�^^�Se�	V�#��X-6�6t���6�55I�C��o�[L�cgq%�[�K������� �֡��.�0��*���ԛ�M���ʑw�Y�[1t ��hS6� S|��w�B0ީ,�!t�x��Nm1��N7�#��T���ze�y�T���X��	h_��:��]Gn-�u	�K�f�Lo$�`�Ĩd1Ol�o�[���5dA�~�y{�E�ܠ��(U���X��ȻK2�p)wl��'�7=�V.�Yi�K���KѤՂyoa$�g�r�+8ڟ-��v���u3U�$]e7���WZ��㰾dΉ��|��
ܳ&H.��KX�>B�l�Ԁ|f���i^��ZI����Ni��]�~�S��}^��جޱP�� 4-�c� ��w6�	B��m�$�1��&4|�h^~�b�Xӏ� s鏫�J�~�J�h��aBD[�~1��kW>�R%�)�>��3�[�"E8:�տ8��龋�=��P��������
�����$��/k��EM�� zu�l#�n����[���35�.��-G�dv��E�	sg��M[�S��i�Z_��i�#Q�z_')+���yz[�Y9B���G+���8]��_�L}Ѫ���n�Wq�I����6�Vڤ���lb)�!*��A�1�~�^�j5�����$����-����w�+�V�[y!�S�э�i��'����}@m(��sE�'UK�Ƚf�jwO��,�F����f˶���9��t;��ܣ2{��^C΃��݉;l5�p,Tܦ /p�F����H���
vD>x ��e$$��zӕ5$��e{��o�ץyD��k����2�n�j���Wrm�'����y�W�q�%X<�9�p�m�תi�N��6���0��-#G�O�+��R���d��A՗�mz[�i6���E�t ��x�E�!�����m�h{���bW^8�g��E(h���E&)x� ���PIH%�y5�����Ј�r��;�hk�#�Χ�*��z� �D��0�@Vu$�����F�Մt�\���Ɠ3�&b,xm r5_��XO��"r/
4�f;���·9��`�+/���2S��hI���o�$�6��#iG���tc��d �ņ�e��'Y�Z]7m�o>p%n�3=�##R"f�p"Fn��A��';�4������AC��@�Fg���~(���i��<v^�v?�d�/}]��(�S@�K��.$�����;OK���¢Y��(&<';���h��Ũ�>'�
�;��o�2�~�Y��ɗ�8FT�`"��	���@B�Y�Z�����M�c5�B��%t�2@��F�~bdb0Bg���)+���5t�B��z��0^X�g���������N�U��FI8�N�q��LQ�k����+��lz��K+S��^��(�������(z����S�pJ(��$G�~�-c��W�9�;M����E����{�NE+�ϱ��z�f+��Y�@#�_��O�f��"�#&a�zf�N�@5a=o\ԎИ6�$��1�/�N��VF��c��H�0� ���e�J�6�����r�A��L��t��$O����H�����ͬ@Y`t��J��1�!����񳰤fh����ր��� ŗ�V���3�����ޤV6�b��|~�Ցu�<dJ�W-}z���=J#Ku�֚��U8����-�U�b>��3�^�;�� ���i�
}*!�����J��Urz��h��j��<�c�G�r򾅶�秚�OfQR�V~�c/�X/��%1���^��CKC�L�=U��38�r���`]�K�ϝ����0�N{{-������u9(��;���r�|��r(��5����K�Z�Ԉ���K-PO�b�ib�#5b�M���n�/�H����!���.�,Wu�[��z6k�|�z��2Y���T*{hΕ{��z�	�EUk7��R4�A�pB�;G6�љ�Ct��9/�v�0��PZ������<��	i��(�~��C	03�I�eDu˰�%Q�}P�<ǭ��#b5�f.�n�H&��F�������*���&�f�9$.gh��[T�x�{60/|�X���26V=ƨ!��O)@` ��C��?������䦴�@��-�l�s̼|
����N쇑���V��<��#3�B�J�����,��>?�XM�r�P9� H�<��u��'|LOG�!��[$"���Z�T�J�A����4�g5�&�u!�?,v�|v@ΰ���8(�����d�n�>�4�g ����u���2g(舦���n�Ȣ��(V��=�H�CGQ}a""P�sYt3��x����W:pH�w���M���5����̂�ƜNA���^�gO�{�j����|E�U8�Ġ�M �|v,��ś#�nb�x5o-ca�l�7�&�M�&Ky�؇��d����um
tS5��2M��vG��J(���,
�"awӂT^��2'�������K�])��I
�SG�N��d��) Ճ�<��K-CϜ�~"���,?-�d�k���NK�'n�����Y�./�rT�<�:|�EK\�,�
B�������y�bdf��������|c�ּyE��̥�jBp�~�����x�1��7�+�iZ �zn@=
�'�C,����g�N��hP��W���A}�Vh�T&~��G���Q�7-�]��?%�?&����t��	40�
v����q��-�ΖV]4y���W}s�W���nܜS�Y,�>4���A�c�+Oun"��.m/ Ӳ�t/�8��f�݈��%L�J�w����`�g6ؾ�$��}�j����@�!da
X��F��2��MT	���-tnyXZ����Y����b��n�`�؅��}��m�c����A��E�*�k�SX��PDSޡ7/`O�y8���B�{��S�b(�5��Y���ag���f�`=b%��n�@0�M0��y��3H�>�._,��  <+�Y�d}�A ��!�̒�D� ��'OZ{��1
¾�Ff�.�
���0�'��චБ���&���Ao��ZQQP��A��&�J���mX�+qs[���[/��Ժ�/<H�Ok���Mo���%."p�B����C�����|�ڂ &�a�,e�Mn\�q�ɼn�u���+E�N��`�XR��������B�!�"�y4��&�f��a�y���ю�Ҕ<#V�������L�!�N ��?˄�1���b2h�ta�IA�B ��0mT�����버�AM�#��H�-	b�6Jo��LG�G�����t���K�cԒ�U��u�gƗ��B�~E�Ŧ�$�5��*Xs�U5	~}�A��E���S�5��1$�B���R(e���t�QGlI|�� �s�\qk��Nb[�p:���cx���8���5:qtxy���������,�ey/I��3�A%x-��U���R���舻�٦:(Q�|i��l�4L`�I��^�&0�S��{IH<�٥��F�G���Q�1������D�ZNu���]����McV4����t��`׈[��!��*�Q���z��"�Hݼ1&8�ӁP�^��	��V��w}�ׇ��ʘw�[�7�W0��٦�S5!��I�|GJ����'i}�g>N�=����d]c���H!3��Ǆ���q2$S��.� c}��R���D�S*��� ��!ˌ�B�!جH���F"����u�AG2sZ�-�Pٗ���'F4�J"�{T�5�,�.��X��R�+PTWf�ѝn","����c��vx�߰�(2����{/8[�u�sQ�XgG�cwdv�ׂ*�E�.��'!��Sɯ5�	�2tZ�2�6^eIj �ŭ�i�`w�z u�z�4�b�B����~�"f�� �4��WrrTt���K���F�� �ФH9�۽I��� ���T�C*�CP0;�� �:"�`��/.��~�ڿ}¢Ǿi���l��wcŝ��.�ՇI��r�3:E<Q��}�V�@}�@�����@��y�FV�g*�)��������]M׈G��-��4�&�Ҩ�9~�0�/��zLR��r���pJ�;��|��s��ofV�6�?Jk�p>�)R4e�i%k>*+����%�$�X{��"�Z!��-{=`�
�ޱ����&]r��;�
�l�)K��� �jG������(3�vUt�@2�T��t�-�]��f�P���d��[��ɰ�����"������t����1�C4�E$�[Ϲ�B��0s�7�VCG	�����`k�(����V_SDO#�[Za���M����@()ª�3d�2��	@J�Xg�ܐJ��ՃV���x�{i�4cy����T[3�P����[~g�T]DLT�w?G02��0��i�D:�����J
��M!6��!v�p�������U��B�놾-J�ni[0hkk�,�$�[;Y�)���K�Oh�^��\+����h󔳦��BO\q�&|��c�
�*���D�����>�t��j/3,3~���&tI=�hj�}4�n�Y�� �S�կW�(��y�M�XԻ�3&���<��S'�n���#�����qۨ&iTw�j>���M�~��`��+^��-7o3w�G=����4ۃ�uQJd�(�L�,��؟_ ?���,F�n�,E��u�2c���K����eD�"�v�ύց��*3�1�SAZr���{���
E�K�gɀ�����z����[�п%x��,�N�3;�~�=��B����]X�d��ߒ���H44T���!@��p��$hSk�G����F���B.+i%�d�Z����fdd�$��m�O�cM�����c�����R$���
���i���ɽe��m�_�$�'�S��no�/d�0��%&��W��[�'�6a�4d&�Z0����q�Gd���:=��㨆w�T^���8�.æ�h���,�w�D�Rt�.��'F��f4+�RwW�B�=O����>]+��b#��`bпY0��4��1T��!k��Bg���swt& Cp�.��1��B�''��I��Z������9+�LH����xI�{G�H�����G)I�� wR~ v*H�$�>���~�l�Fi>�Ǫ3��SǺ��I��eۃ���� �wg���X�Z��nܰ�=,G��$�b����D66�۝�r��,^��%A���e�W����C�*�W���5.�78
�Ϸ�����nC�b�{��W�}�>�����A�Q٨A ��������i԰G#*�K�*�Ң�@Ч��-:����9HP\����L�ac�jSk���e���΅R��X�m|�"�lB&-mΦ�8���4S%��b�x����S����D[���� +�oj8�b�Qc-!��Ɋ�E�C}�e���Ā�9��V���G1�S���]�c���|(���Ĉ1���g�5w�;�0^�|=^�L�-'�Cg��n~�6y�������i�����v?#	�eI��0�$F].Q2@5w��Id�s�K�L"��|�=M�3�����6�77�����y`V��.2PE�c=�k�Ѡ��T��H*��]��]H�R�[O���݅��.3A�LuR{��RoX�B4rp�+N�a�I�E��~���ʋ�ݣ,�6��y�ۑ�G�	�HiqK3�E
�}g�_�x�rLB��y�If��5bb]N�e��i�������2���d�F�����K�p%��J�Kʴ��z�N�@���j��x��5�ޚ�b�qC=�~��Γ�u�K�N�r�Vq���U�Ţ���۠��N@�:jw!�	� w���#���E�wr�З@9���%�{�kA�.�݇/kx���(=ԩ!��+r)�{ѱ0L5�ý=�	踍~���재�z���a�${٪�b1"0���`�����lε�;C&���#��F0��8�@a����ː�>������5�U��Do�$��BhI3�-��>Θ⦰�G�]�@rmT�n�f9o���!g�L���I�S�fd�`u��ZN&u",�Ov�O|(A'r��KL^g,ӨW��/���D#E���K ��#�F��Y�|�<�f�,���j-�~��Ue��@���ko�դ��<�����q�����<���H(�v����g�@FJ}_��Y}đ-�टT=�Y�N���u��t+��3c�?��Z�^��{�U��'8������0�p�`b��Ǵ�N�y�^��8�F):�cby*��G��s"սn�)��<�٣��$�1��\�-J�+��b\��ڣ�.׷\ �@\6xV��/w�nR��>�.�pY��X�#H}a�|���w�YC3�S=�$_�I�{��!���H ZZ}�>������$�l7�6jD��s,{���7�N?+��d��W?���*��ĕ��ʯ��1W�%�dêҰ%��l��@�I&����/G��w'Yk0t��4�%�l���5��m{�<p�$ӈ(���3��
jg�u"AO�]�E㿻�ԝ����!{���O�Z�mfrٚ�O��R��Κ����3v>\ϺW%�x�J^��0���,������΀����t^vW��(
�7ʆ}�N���g�����*�]/�Qq�1�k���]B��a��@F�&U�u'�͠�ӻ;uǫ�LZ�Y>
���ل
8�.?WTi����k��k�	�uY���� �W#`H��'5�!�z��XRҫtzBWD��)M̺��B�o�$4���`�:]bCs�k2��vp�ߙ6�*�vL�LRy@�mS��,#*l��z�@��]�Ŗ�p1=���j��Ych���ݲ1����w�������b�e�^u.idǇ�����6Zk��2����%
�)��+G�R��$*җ�*�ҽ��������.�5����_�����>fd3:f��hT\y/���<�a� ���t�p�Y�1�Mq��Ⱥ|�q�R�e��E�Z����-!�E�S�+��):������L�r�A��	;�E���#w6�F_辚W{���;�m�<��1?)�K: ��	U_�Pn=��&��j�L�l�
 �Y:�R������#$L�3J�R'~�~o�3�פ���~�.;8�~Ǻ��Ԅ_3��!�6�65��&�����Aq�G��4R�=���;���(���{␲��}Ƈj�Lݕ�M]���2erpd��W�ʤ)�����'�|>��,˭B���e�3�1b!����B�<��Tn����b��&��|����b�r����^zZ��q��w� �)�٣��*�Zѿ���k1�VX&> t��
��MI�D���n	�͙�M���>�;�b�8	17��Nn���4ү����(�}�V���8�/�.|�q�i�ꐠ����&6c�6�q����Q���f����墼m�ǳ��5��vE���q(�`����m�5q]:^�r���c2��k>V��[{�#>�Ij���D$��/j>5Ӂ�!�H��~̙���i)É��e�`�����Z��vK�R뿫�`���<�P�����<�P|PY'�ׯP�vF>#hS@�(O��޳~&+a�F�*��ѹd�$wj��;�L���F���b�~q��Ύ��Q�,|mG[���g���<��^%���2�&lh����$y�aZ�l�G:\IJq.s⨃�߃3�)%�2�n8u	�P�o�;���_T�h�pG�Xv�i#���W��D�2+k�dJ�Lt3�A@�E=."��sF�E���������e�yo�m�n.��v�a�Qsr�[�i�d��Uy��`�c��+K�lF��~\�:E��?;U�Z�s�4���k�^q�w����3��*��כ4^�].��L؅E=������t�H�L���F��R����|ǎ�5�*^�di���j���Љ���~M!�$��>�#���(�>ġAs�,��|h(�I�2H�m�9��r̆ӑ�Ԣ��h2����]��ZN�Q>oB�B������޷�
��2��d_}��F=�)�힍�������T��� ?�-͑}mU-�RsӶ����+f����o5n�K�d�[��S�!���y�X�I��"�����@�FGψ3}�*u��lV��t��TR	��/r-Nuc��Td�w�/xD���b�PR*���*o(���)4z_}dɄ�/'Y[$��!���: l�0�%�+������&��I�b� jα>?��?�{9M�e�c�b��?R��b;���o��[��V�D&�:p>Bn�����5��FY�z�:?����.���B����è�'�zR��x�t Hv�hr��P1��uf�i{��߹f���6���d��2�ĵ����r��):�h��b����_����Z5[�^�0mmw�lH,Pp�
?�\\Z����i[��\n�
��G�@���Nw���K9C;8�pA�vՔK��6��97¬��҅�n�eF��C��K�H��Z�夎��;��<��+`9�K�PQ;49�na�k0����Y|�HL�X��j90����%��
�����N���ˡ4?��I	ڥc�@�A9�e͵�L�FVMXj��i�JhZ����[��;'�������0Q����ҙn��	f�i����A���"�)Y��u�~r�=8zٞ��T�(z�:�?�r��I���bT������r�@4�ڸؙ�!������"H�/&����9=�:P�����;dĚo�ӕ��u�|��ˮΨ�_nK)�+�̯��������7�܇�Ic�������@T�;=o=�M�����_dp�\o_~�(�Y�+8;���Q��)�wZ�-��x���Xf��=��s{�6$}��W�6�q�U�� ����3{������#�І< v|�I���JPZ *���9ETi�ܵ���+�g�����������OO��.ys�[Ъd����7zLy!'))��������X���6�q��H'�Zw7B���]�K�n΁�R@̎�EǡS�����u"�X�|��p�O����N�E>���J�d��i��t��%���0���8�k�/�G���K��5Ao���	*���>M�\y����i��Z���a��`�~��`O��^�{�Lw ���,�]=]�D�軎�{���W�������Q� �[��n�l��t�L��R��/�mf�nJڝ��M?����/Fԥ��r:�ji���9�X,�Xr������Y�Vx\���o�FB�;�(��a��2B��T�o��	u]ydt��?Ql6��X+z-�(�yNvv�6�L���,~"ĉ(�1��J8�F��GFZىl2����7�,�4>��[[��$�ٹ������Eg܅&�XJe2�k0H!H�}���A�UO	n��~ �����ta�'&h{ox��x�k�K*Ϣ�Zm�a���+%%^����K菑D�p�B����y�!�_s�����X��_��&Pt����A%��0I���:�O����C��cR�[�`���(���"v�d3M�C3J�g'@䙭I���A�r�/��B�b��~���֯� S]�ե����&|9�26��b"��e-nw���{�~��G�mKt$}�����)cf9����.Bx}�K�A��,#b�nm��j�8����ɳ�Ad��S�1�`���Ш[[�吴��ؓ����
 %�2��Dd�,`*��1��s�xpv"?�Պv�oAB;YV�������<΄�����'�
����p�b�W���H���^#~h3:�V�;�����"]^G��ٺ��k��k�q�4 }��߷�(��Ѽܥ�П��nH#a֋�l��(��b|�؟�����Kz�i"��ȣ�s��ym����S���M$��Kw���`e��@@�ñX�{-��|b�~�8�U8��k�=�������:�/,`P�g�,]bE�du1��z�j������fNS+Z���ۗ�vNS{�5�_XC?K�8o��Y����m������
�J|څ�_v��cy�X볝��ANTP��0va��p(h���1&�w�鋎��)�>^t!Tm�OQ7?���7���MX�}�!�L�� �+%�,���j�e\z�2Ю�xƖ�� �n!e��pgٹ�sfx*����iko�N�� n�1@���+~�VQbEw��j�-<b� ��l�,H{�����Wi�����ԕQW�w������l��mܯ�6`��� �+t���Z37))��㫫�d�kxǼo���e����m{	�_�?$�S���ĬG
E�e�������C:���=zI��E�	V�Gy��D#�t���a�д�9a�W�cw=_�HD��@q��-�{c����ߺ]�p���}���e�R 6�� kW����ԧ<b��L�M��UMjMY�T��x�fe�J��pӯA ܾB������S�+��}~9����-H	���XDq,F&�m~�����%/��5����՞p Nk��r�����r7�`u\y��w1ى2����vy/>��%�Lh$kb��O/9���9Uz��w�߅3|��I�v#�A��I��<K�/Wl
��v�_N83]�Q�� i�U`[]'���0�9|���F�ç��f�h����_�b$�d^�*��ԇ���ԁ
۟{2T�l�#��4(0�БZ91�ޠӥv�Q��u
�n�}g&?�N^�K�+ulYu
�]D�3���a^Q���1xO�[8Y�Mt� ���'5ן �O��i�����i��7�����Ϋ���kقX>|�Z֚Z�\��"��rV�	��z*�D)5Ы�c��rk">.��{6y!��t8��x�S�Z,��]d�4" K;$�����I~��Kx��#?���A������>���*�
���H&��Z��yӋ�Gl�T�\�4��8w|-�^RR��ʝ�w���iåՀ�RZ�PZJ*�z`�H��'�,�ńM�EC��S��v���V�ը��� ҄���;���~�W���L�7�/;b��m��D[�=�^ӻ/�Ѫ�A۬y�褍ϭx|��X!��7Cb���O� q� �s�V+��փ�!��ɍዺ� 
�>��
)���k�=�3���V��H��f��4o�9���}5�=j�_���]N.�����':H2��2Qo������^��3;�y���o{�	�?�X���[u�s��9�k=A=���K�«�<(d��Ǩ���f��l�g��s3{\~v�0�cԸ̷�j�7�����s�S�&xVs����k�$g�L���Ĵ�D�.P�&�
ᾕڅ�p�'	 �r���x�ZCk�d������)%K�Y��]96����Kzeo4AQ�G�n�վ ���)Q�24�4���A�p���ʥš�!���h;��~�������Pt�L����3Z`_�)�n�$�$.�(��N�O�پw�9k4�>���	-��(�WcJ�����l	L�Roˏ/!:��瓓]��ZI�Рt�&q������#�X+����`��lWq��f�OzhՎ&���y"1�'�D�·�Q p_����!a�쏷�a��^)��4�|����ʚ�<l�`o�"G��T�:@T2ϩp4e�?�q̂hOJ�4�����	N�[1.�V�� ���6�Z���=%[`��%����e^��[p�!Xg�~�X�0��z�0��΁lbކ�(��	-3���K��jN�i�06��н�39 ��` mLnVt��������ԥ����%%�%\���R:�ڑ�<�;��u�3�X�u�sW���b�d}�wi�i�x{cy2�ӗ��'\Y�����Qhr}��x�3�gۖ'I)��P�bIϟ�3;������K���ù�=;��6#��G�k��PJ�:�/��j����и��lwz*�a�}o�'�v�)ʼ���/e-�h�/v��1!�d2���ёj���|��_~"_�8҆%��A� �s�Z�4�����Est`�w#*����y�<,'r�wd�/�H�Շ��Ek���?p����_����}Ʊ4ݐ����=��~��@�M�1��z�.I	�U>;��ݮ0�Bڞ_��Co������5,�ͩV����3�r�k�mQ2S��u�obF�W��S�'�"N��H
͗IQ�:1���?An�"���l����Q��¨��R
tS �@�2�CP��nC�A�&u���m*��7��=o0�>��b���.$g��E)� �����8��!$���;#�����P�<#ŭ;r�Ұ_��F�m[u��]Q�M��ۨV�����U���A˯1�3����ٶO��l���'��B����k���=�R3�]#���n�T@��]�c���sa-Ćy�K��MJ-gN��ρ,�g1y��<5�M���M[q��k��L�q�\�G��:�����U9&�(�k7�{���X�_�Z�r4Oh��;2t�z�` u[���A�c#����GN�����Re�z�_�o���s^1�PI<)���2���	D�yc�D/��i�5U������2��C��9�m�s:���ʰ����(CЦ�����z;Q��6�|�x�f��>l�_����
8&����"�緮 �0!��`�/�G��Xf�{��u`�֊vB������ ��TX)Ta;�x֌!�r���	�2O%ի�c�������i=i�~ak������Y�_�bu��W8(\C��Ò"5�nIB8� h;u��_�D��2�9����`�V/���ȅ��4�0�:)-K	��QK~�7^� .�E'�r���P�/�	�;��,4%C���R�IS��A�]�]%�n΃�պ}�mXsNm��"�ӣV)��;/�,nw�ɕ��f�����"!J_)mf����>v1��|��X�����	�,�_�o�m�Sj|EA�O8]OJ��m��܎�}�>Y3Ѓ�I���U��,�y���d�o?�w&�a���s�;ˇ���-k�;��ӡ����eD�+:2t?�,}����V�v6�5�����̙��r���S�9���h�6������Y�zH���q0��E5V���	MWa�\�n�$��b�t�$�"z�m�GdBN
�gG/T�Ù�O(�b3�Sˤ ԛ�*���&4ia8kH������ȧ�=�Hgv�y�h9�W�R�<E��)��t<�c�K3֪�W��uʶ�O�Ui�X$&~{�#�p��ߨ0������5b�){-�~l�,�M,Ks`�B����補V&=�{�>!t3�al�}�L�\ˏ�bM$3��A�w�/笼�NL��ު ��Fj1���b��&��n�f��^:�+���'p�f�����u�	����d�U�ўK68�Š��������ͦג
Q儾�Bj�,�l�Ns�7�$�@@�Ҟ�#�l�H1�c��P�O?��#X2|�@-�<І�<ΐ\���`�F�B��/�E�dE�d���#0I��M��&X�a I\�m�ɗ��k؜yS��i�j�unn���;�"��8���vu&&�-�avy�9�O��蛈�AT6���d�3�Вܬ3F�W�8�M۱g�/�F��I�І�[�^(!H��y�g�(�k�e��Ү�l�W[�eLu F����ߒ=��x�莳w�Z�ؐ�Y�dӁH@���)`s5r�?�Y#1y����k?^.U:@��GA�a�y���'�O�*<T�� r�R�,�TR&ë�ز���041�Z�H���=9H���j\�lN���b����2���-�d.��:'o`R��Gc�#�d���Ɔ���*��鍇�c�Dݿ�=��nz�5K�Vؒ#1�6�����ķ��Cl_�KD��r)G5�)L�#Gf����-�Ҩ����;�	�?UHG��zr9W����� ��ܒ@fy�b`��pp={'���D1�i����*�yc���ׅ��#zF��'��TG{*Z���E�x>!$�N���������@��O���z�t$��<����}(�L��T`-z,�Ed�k�d?C��0�x���¬u�b�7'��M����Az�YZcT(H=�m~J�#��i�]o���r<�)R�O�`�V����6��Z��������N�`I��@�u�ŭ<q���8� ��3�8s���*|J��&�@#��h@2Z����W&���5s��Hٓv�v(Nk�/?�A�Sҁ�7�6C��g3�x,*z���4ݡ8w��)����6�)^{�����G-���?��>�q9M�U�fJ��H!x��}����V�|��<�x�d���%��.D��������+�54f�BIK~sP~s�mhdמs="7S�d=�3}�1�:�0�U��$PN⾼�G�u���1Mþ�Ό+qm�ηsfkMmu�ǒ���_O���n��E�D���Yd4�G��	���Q�?�o<(���W=�{�4���xCS�_U	���-�_W��y��)�yc�m�%�}�x�-X���o�y�E �G�&������:�	�e���^=�)��\�v��V�����q�3��V�-��}K�-����,�&%�j~ܭro��ƨ����V��z�[/1*M1�A}�şI��+-�;�k����ԣ�ns}��fJ��b�5Wf����wF�������6�[L��J�����M�H�lF>KE�6 ^���{�����H���L7.Ԋb3�18R��������\.zΚCtͥ�	K���I��*P:Py���a���#l����:9�����8V�Vodh�I��H��nx�׬ ����������4#�DHE �WUMZiY �8�`�!Q
l�/�=����]�:'#C*S]cpuT��^�&ԗ��>z��Tg���}�ڃ��l
�)b�M�%�'4CX¬�G� ��\I�]/�Ҟ2>��^�ߺ9��'���(���$[-W���Z�fs��K�!�M&6��Sbru�~�W����W�� �?rF�j�I%�C\!'��r�f6�lJP.�NE����<E�[&�������j��K�n��O8�t����S�Х��uB�Qgה��!�l4���d0����rA��ūY[�IK�A��bͫu�������
͏�پ�i��{#�s��Qf <��i 񘻆��e���<�����h\p�lU럴SӹO>��265��`�*��8_6`Ц�9�q���t�7nT�M�����NWH�כ��}�L\��wEg��T��?�VK5�/�6$�<��1Q���g���8��.��e,,%7�Zо]�!��m���4n��������9���p܊_���o�q�EM�C�,00�;��)Nu�߭��ug&(JڏvW�F��'�h<�i�9�������<���\�
�-�����{k�� T�D�e����@��t
Nd�p�X��e�Դ�-p�6��D���v06��+<��^?��R,�:��i��m��/һ�-U��Y�vM��N���ZL{�4 ��*O$S7}py��rI4�lC�-��<�'{q[?���|�;0�p��u+���Ez�[�� �A���z���tb"�]]'ɛ]���>�h�Z$�7+��2��sKۈhR-���o%N�%�j�H���,��m4
�g����İ�	��:�y�P8\T0Qu���T@VNձ���`G�Que��GVW��w�id�yt��Z�����֙>1�Ke����!�V�Z�S	F��j(c��Ԯ�-�7!~s���B�XH�sOh��H�s�ޔGL�-<	\�~F�*����w��`�m!��d�WB���ʓI����dq�����mi�f	�hq� 	%��9�!n+�Y��T��4�u�F0H�e/CܢL9�*��X�3	����<0nߎ� �{�ߵO�w��BRU@⸃�W�e�xg��ȣ1���κ4�k��'�m�}Y�el.�/%��>��0w��he�2�$=�/�^�����!�!�2)����܎ؠ��F�Q��C��/�/f�\G��i�)���S3☭����3Gy�(GU�����}�)-�"E�J^�ݩq�|r��@� 5|�׫05��T��V��f��p�0z����6#l�&4S�L}��)d�t��I���`���C��7�P�|��؋<���(KrEڤ�4�Nb3A�O\�|�Iz,RF"��3�Ed]g�Y��׹%�i/M	����2Dfm� �;d���@ϰd��R��1�xzf3B?<.r���zk��bv�!-���9�Qܬ�Ş��͕���~}z�eU��P�q��u�Ծriu���� _ ��2��4"�1{)�*]{�h��&m��U}v���i���`�F�~,����
��@�ℋ5�SΑ\�}!�9G*zO�����R�k�."�RJ2�	)� ��ɕ0.�¢���OO*�.�i���1���rk��� �;.���OyN�P�������Mh<B��u_٘]nnb����L�&�S�C�搻0�Bi��6�)�����,�Y ��rd��'�2@� ��/h� .N/*7Y��j~⑋f��:k�_�=1U������Bqa�_nz�8���Q�pzt�9*�9f���n��]w�S�}-���&?Bk�%FsN����?[�Y�z]�(bnhU���d��C�j�8�^�R�p���w�=I������z�M�J&F���nܽr���3��p,}���u�)�w�>�N���*`�MT�@�^&�S�����HX<�=]��h)���(l�@J�2s�+�+�S�4��v�Xg�",���Iؙ�<8]�.����Q	�G>'a��Hv���?�d>�Q��O����4��q��$�5�?�� %���K�<+x�s��ͷ�P�
���j%Ur$剽��a�ɬ'�0,Z
�j_��y�����yr�Yko���2�X�s��9F�2�>@8�!=O�N�u�� ����0K��fL2�;�U�~6�OV��Y�mb~�Xx���̈́�T����������Q����;���ªX�y���j:�;*nl���w�d�@.@\�DdX�3�9KU?�t�&=�ށ�uL�}�(yܣ�
�c( �F�-��M�v'"����U�Ơ�xà�}�7�=�z�v��Y,N��gM4}�	�9U��.�2Π�dA)#S���U��̱=��fP�� ��4E�f�t�[̞��5�����5�|����iH��/ �:�(P0eG��h��N��-��SY�[X����j��7~�x���ં����~���!i�V+U���@�T���(ˁ*�G���k>���#o=t���%��%w3䕳<�Of�K�5�+z;��t��(����ϻn����0Y��6�/��ȹp��咾A��nl�V-��W���)/G��,T����: ���F&�����ȕu���hPR����=���ҿB���/���n�܀d�m�'E���a�R��N?�x���
�5#��t�.u.�a=/�U������c3�^�W��_��j#���'b�D�nt#���*�"Hr	DQ7B]L�Qf�SS��s$:9Cxw��XNbZ��)����j�m��^ ?h�a�n�_b�rK��;k�>��!!�Ӻd�����iA]���;n��i��r���K��T�yi�R�\�:?���3���0��BTV��Ա����yn��~�9�ыK�>tƣ��z hev��9]Z�G����YC
P���nJ&�̧��F�𕏍��b���@��T^ܠ���p���tP9ŉ
G6\O8t[���H�U:�e�z��4�`��������������2eR�fDW|�|[ϻ��D8.���ݚ*.�s|I!�>�|60��H���vojk�/Mdwg�{�*�Yte6�!Z�
:�e�9����ᾃH[G�RYrݷ8�y�����z��B���PJ����u߻����s1�Z�ZD����R�c�m�������a;IBy&C�ͅQ�x�$ףY��Ĩv�|P�+�Y��T�Q�Dpz4��Πtr64-]�M�.�V��"���:��1�� �@P����O����(�/�O�![�[k�@�c�w9L\�8"e��̾r�`.�,Y�>v�?QZ�S9�P���H���-n0@��}�R�!�7s�/���e��X����a'��!���]�E�?�ΐ���$RYr���Y%ɮ�{�jŒ�.��E a��1y������!������gs.�߮ȫ�r�],�$c�]*��˔��h_���%����թN����i�}[`����i\���a~Z������ ����N����1�qa�9��@6��e׀ĥ�ߏ!P���TҹW�S��`����#M|{�$�C�iɜ��3�#�&b�;�w�OѢSx9[����*,d�c�ث�����M�=�K��o'n�� � o4�{��V8>�Z4S��O�� Pr��ޙ�(���j�op30�3�lλ���G��Ѕ�����+/om����`3z���4٬b�*�@s�J���n ��Wazn��!�8�xR����"S�b����G (;m�n��{H�ѵ�\M>���~���mؚ����eG��뾭�&N�~q��>�2HɃn�"��p����Q�uV8��Z	�9ڤ��#�8p����Yi�^Br��;��ޗ�
��m�g썬o�waS���l|��+�np�������e�x`i�������*w�,��:�o�y��{�����&��yp3
^��ݯ�Nv�m(���*f*lҚ�f��.�b�^��l���I3v�~��a����-�*ZlT��9
�}^b�g`�Ǔ���(�,�/e����艚l�i�gEl�fث��CE$~X)������[�L�ye"-c8����M�ěr`g�j!�ǟ�	�cf����.�Q�,����}�av�-7V��a&B�nM�^�_�<v�D���u^b�7	�Ж�zơ��c1�M	,�;�O[S��\��c򺥩��S�)+#��;ΑGp���|]ogJ�(X0R�ۤDK^��~�����q���{Yʇ�-!'Ȉ�'�$��=����A�_��_��������^��z�j5��B79� ��4���1�(ؤ�=x;�t��b9�i?�d�C�q	c�!�2X�'7�_���zs^�\��l4f�X���`e�龿�ʤq���������TM�r]�+t�/����:��~7۟R^�н{@v��>��m]�aK�w�1�4�r7�f�]�1����Ǿ'^ �eȿk��MЏc7�f�hRn�*t��NC��4����z���1O�ϲ��\bA->���H�ߜ�>���&�c9~J}%���2ܷ�7I���t�h[.�C^R�5�wJ'lI|H��X� �;cƢ���A�,Y*	��&wΜ�/��U��3��Y�����/�-Z�rJo-���t�rVUW�ck�[JL��@��@�6�rB�2�B�A�\;�����t�.��"�����艩o��X�@��$f��?�fb�St�	�3�ifm�I�ܸB �X������Uaw��#a�S>�`��$>�1Q�X��UR�?lZ�/6T��U� /h^6'{j��ۢIfJrY���bܺ�q�\$�N1�L�~�Ft#T��}]��׆�h�}}�0�_�O�v#0z�yO�:CJC`����5���
��mʥD(D������ǝ��o�24g<��Ͳ���[^��F�N^or��� G$����!�If�,%|:���g�2����tg<����&�Pw���9�l��
ԛ��*��s��lO}�X��+lN��"{P��˱C�\�;�B��d�Ƈ|q,T�����0�G��B��8RW�[���R�������K����H��ͶT''����C���)����
����I�w/��8ڢB���n��l�B�kS���n%E�t�0pY�ɜe��8�eU>/��%�"��9�R6�"���p't�H	����L!Ǎ���4��3�ec�(�?T�mV�y���CXV�Zݿ��@�s��>n����;<�F%�V·���1��}\���GF|v0�\iX?��t@�Ԧء U�$���,���CYӶ���-t�"�v����@7����_�+g�q�(l�.�{�A~s^����������s��E��6\B��I96|R�^"Gu
1P-ъ��!�D�@���l�4@SI̖�}.�k�ɹ��N���C�em+.k���Qk�Xoң���"v;zGzM�IE���pH1B�M�w2�>����#~2��������3�x5���	7������y�A����4�R��Zg!��V�Uă�1��٦3<ZsaW.�~�/W�	����%��j�7����T��e����M�u)�g;���7�:f���Ja��jFl����v���u��y"Z!D�x�Ĳ���-r����}*��3�N�Cx7'eV�Xs��xh"~�����RȽНU����i]kO��Vؔ=���
p�uI��{=裰p#|�c8 I��*�qF����\~�dQv��Y~_t�[ˑ�KYL�$����ي��B�� >���-2�چ^��қ�P��+�<�j�e�m�CJ��'��G�q3w����V��B"�"3��0����j$�G`�2�Jt|V���Гs�����k�㴘�6�h[�p�'MpCVPP�k�T���!}�ɊHz� @&�}Oc���B!"������6��$aY���n��f m�D~�m@o%���P�o���;EC�y[ �,���ٞ8z�&�	1s��0��~`,��ɲ��rP���iDcW6��� �*�4�n��=y��^ʹX����j��#&1f����
�T��ɛ�2�w-�����>%���/xP�:I�� ���������h_�Y�xLƷ*���%kY8�pu�k�#�	_۽���c�>�!v�{34��F�U��pj-(ݰ��ύV$��~�to)�d�Ѐ�>�e��7K���{	[1�%s����oi�>]���O�`��$�@��
��w��3�wy�&!B�B��.;��J��$N�i;�^����Tà)#"��y!�jeM�ou;&���|��u*q�C&i2����=n���T@Q����p�$���ѹ*(�|�"��#A�Ą�a������u+��U�@�A�-{胺s�Xqb9�����7�CtA��-l�TR��9a�ڐ�䦍��m�g�}Z'i���ن�k���\�IC��-zw;]�a˦�|��%@/��r��bHű��Q|��vN��ONUZ>�t�2���v��G��j�O�;4s>T�� ��S��(	8��
��S�0@)���WK� x-�ewi���+/��宬&��H��k�"з��u��R�W�Z�A��z�7��4�3�<-o���2wjfI�"xޣ��x/�T���!�|��F��˅!�<'}�7�6�m�@�5��g7�����ݤh���#�ӣT�Q�@���}��(��ݒ�hEđN�=�ʙ�/Eۑ��[P�ǴO��P�3���Q}N4=8H������>齾+�2J�*q�����B��9�t�,��5�|�O��OS�b$�6VHq���y��j�%$5٦hV������i�E����T��R�PL\	���1�G�Z.�4O�a�F��M�![-��GӋ���:z�ǐ��x�� ��;�{!q86����rKI},(�?k�o֝�k� �<JhC�D}��ߡ^��N���c�KN4��1N4� l��`Xy�0`i���J�=�#PF��)�PB�J�!?�"Do��j���m�O�	O�Zp�N{��-��g^�S�hG5����V�`�p��"����C(�J [�jI�B�q��<�_Ȫ�	(������QO,K��'�^�Y��7R��dZ7xNt��.׷���v7������ס�ܼ�v�f���-�QDpw����b��h��h7ꓞN�tfh[���ԃ�Ӹ�'�?��ƉA��G�P!�_[UN�d%*:s��	��lş���u�D��OXB�.fFD��0�s�C���t􁹋)	��:3�_��?�	���<p������R�|�B�1��Un!�"�9:a�)P^_��ve��I��+`i9,�Gtռ�L�����\�Bȁxoy���-����Y���f���=��:�G�[wK�����x�8l�	��7T���	?em�<��U,�]�,�&���}=T��Vw����.�bÓ]�ݖ3�,�LBA{)�G���fkL<��,�Gy:6x�sh'�2���c�!�E��{���(L�(�b,�������t���E�%71R]��'�K�≐v�?�ſ|��6��b���@L)V>oL�,�Ε��O>�������V[һA`�a-{��o�u+Sj20N?���#A�N��M�
��<𻹝��A�`^�7C�$�	��5��z���u�h%�fu��|al�"�5�m$HX�-t �8L��$�� d+��p��2�}_.J[�$+���$A�3�A���5;��(n�h�Y� J�R^���s&���8�"'	�`�$���R��y�O}��4[\�Y��� +C"�糾� �ƶ_��=���V;���!~f�f�Kc����giR��ͨ�s�7dy�Ե|�;
���щ��h;w��_���f�
H�C#z��=jB5_E�M_�A���%�z��_� SE�9�ݓ��uޕ7	���:��L��^{^���]�Y6_��h�_M���'�^f Ci䗲[H!3���w[�׌���_'�E�� J��z�K3W6!���ܻ<�K�`O��Q�d����e� �K89��i�Tc٢`�Y&�%'��B��$�NMwk�������`���	�R,�Zx\�``��!6��۹�a"��,�_�'(_r�������F�5���z�~�|IOmDȊ+��dؽ�ro�IN��P�?f��2Yۢ��X�n�G $�uo/<�|�kpM�d�/�Ie��LB�6=��q�%�	o��.a��+Pԋ&�<曱*��!?�,ÔGz���\X� ȴ����)JO�k~)E����frl���5�"	���Ր>�L �����1xɁ�xy�`��>y`s]x��'�j+J���E��t_�J���`e-!|å �~*�0��B���= ����ƣ�ڽ�^�ͪ�ʞ�t�6���7j%ߟ��5�s�L8�l��)$ў� FZT�:�Ft>��Vi�lѲm��{�d����&����Фe���`Y�k;k�&�4��ewf[�g��O֡��S�.�f�c<a�8�Z���b�jDco�c!IA�n�����=����q�C��9�j�k�W���B�i�Ű�&{t����N�$r���p2O�S��P�	W���<�������g��w�����(>wa'�=u���m*֋�?��s&�Q�R<'~��&�:]#��];D���KX�d}�Vj'�����S5�OL�?"�B%���7�vIx�P��پ���]�����R���*�|&=�٣���Z��d�ʖ�A9	��$�c���9Z�	�w��B�D�P�=�"��/���C5����I��^��E�&g��r��5�Č��� ��.��Oހ[W�T�R��5+~mӧ�]���ڒ]/P�NP�S=��Ym�⺅�(Sy�<��3g�>�yL�G�;db綒h����t�[�����\5�����`U���� lS1 3\�x���+�!^Z!�̫f�X�8y1��Q��u�3P��BU����fF����:K��|?� (~/�?���/wQژ7�D�u�F�z����N�d.
P��MOG�&9]�^WW�@+(� W0����]�[6Rw�9�|����Td%
�W�ؔԀ����Ə���ҴH+��/�}i`yex��	ϐ긒�����֯�CA�_�q�d35����#�Haj�v��'Һ�.<R��Q�2A]%L�_��D�5$��!�z���2\V����kNB�ӏ����<'=�N�.n��L~{q�B�����*���#��I�z����&Xjϧ�ҍÌ���d�xi\3("�Z��@ێ�З��?p���
%�6q܉SW%2���W��e�� �ϛElh���R]c^�@�@g��丒y} 0��YWsK��f�T�6�>5��^����3B���`�n�Tp����!�mS���0��k�g{���� �P ���۩#����8ά�|�Z�
�뙝�����%�r��h�J�7@�rVP��@��<�R��1Ɍ��[���:@���q��kڽ}ٝa���#�Q6���nC6��6:շ������/��Yl�����I�ڜ0uS��Yiw�.<�dIwr�0�dSs���l
D��Ѣ>效�`ܕ�X}I%ɱe:z�AS��j�=�"֝���j��3Y+�^J9�u��?���<e�~v!B���e����lUi4h0�W���z�p����F9I�H����&���!(�~IT����f�X1(��b������jF�f]�D��M�Vad�>Oz�4<5����Z3�$������H	B�����w5S����y��IJ��2��*�bG8���i%� �0�M#�R��B;'n%V�#��:����������tl�uC�]M����|Ӕ��K�_ǘ��p7I�&�|}���ju�߸S�~>e� ��ݪtG&�q�6&6��7�s3�?�ZI�N�n�6��l�Į� �U|�jhA��v�H|�GG%f��:�a��E�.�W�(1o�������d�/���'��:[Oq����N+�sE��0�:a���*��WI�T
�`�z�����95�H�E����GaW�L~@;� �<���+�&+�vx�m=|��H�-+Q�����+qͷ�(S�ל��}��<�k<C!jT&ѽIl������Z�4&��q]���j�V_'��B�Z&�ȂE��b
 ^� ���;[��[˭�rQ*��K��x�̼��Fw<�9]���Ĭ��ˉ4��q�����V-xj�Dr�78�-5���Z��L���=����T'yjne�y���"���fƵ<��^�5����u��#��4�4a�47�C�b=��Ы0g��H�;O��|wxn���[j�rƂL���F�{<[!$�%s�q�k�kc�n���evt��4�Z�>=�JR\�O='���&o�n����${�u�SG��ВF��� �&Mt�ʀ�i��2ᬘ�S(������^��[|��
��|��o�
-����O	��&�s�Kխ�G}�%ϕݨ�	�����n��jB���3L�%��@1���|�1���x3fc-2��K��څ���!��iwk�~㼞_��ć�dީ�2I&SM�79��6��D�u������=+�'��s"���`ؙ*��=��LD��'gB?�CZ��)�R�'sz,L�2%���y���c^���X���k;���KR)�r��y0w��:�pבB]Q�9bzm*2�
�89��P��<��g|(�� �$~�p �ݢ���n?u�(x�����Af�d�hc2)�Jz!=n&�N�/�2J��f����OK� S��9��>~���)K����H��M�A��lF�sa��<k̓Iꯝ�!oU�����_4���0�OC?,nq�/�b���&���":��,p��bFD�a�.M���	Pn�c/cv������<���,�,$�Z�s��X�ao�7"<K�jB����T�n/�*���lç��J���|�+\�a�;�)�i%�����W��.��sU����/�Ӻ�]��Q�ɂ�scϭA^4��*N�:�lmWn��N�F���zTӆn����H;�^�����r(QjZ+���
�MgʟG�cý����M��&4#^>�ifJ�r1߯���]7�lW}���q)��j�"��3�Gҷ���.bw��[����W{��i�|F�$� M����66s�[&կ��-���W,:H�J*�8�8�N�� ����3�ŀD��>:p��F5A��7]�Ňt9��)/dC5Td�x�6tB>��FI$T��@��vаĥ{2��,0k*�ʜck�U<K�?���{<C6���ü�������s=^7�Y�3��i��.3�k�v��ƙcr��Fg��ʺ�o��ΰo����S��zK8yX���7��c�������rB��1�h�"���P��Ćp�I�ǷK^���(q�B���']�֬�<��1�]/M�r4��;�$9u�h��*`��I��Kk{!�y���*��
�z��9��B�#��ߩP�peW4n�9e���n,è>�ξ�ݫ'�mE��:���Q�ji)�P�܇�02�jK��l���6b(�]�����Y�^�8��];����N�*C]t��%��a�9o�]�y�z�s4�8|#��jsUx���Y�q8�����p���/��E,�KYQp���=s{�v�%��V��NR̍t����['ԃZ�˨�DB�T�.[���ki�fY�c��Ww��sd�N~CU�	�Q<�,��l��)��'���{C%>���g��?��IҌ��j��h��I���BC���vw$/֕1��=~���+�joe�Vgr�)4`w���aW'A֞�a� ��-g1Asmb8Q$S�ִP2Y?k���, 	��`�C2�=1<��BQ���A�l9-@�����c��a�%Q�G��� �(��9K�u���2�|݆�]��Vޮ�x�J�$7��Xx"��ޙ\��ݒ��xԔNB�D��K0�ތ���'Թ��/#z���V���/�&�q�n����kdQ�W�N�;��G�)�[�������+^�"ܯD�j#M_�e*[ܪ���b9��R��l$�P��5��Q�?1�����p�*Nͧ�H֤}=�^�����5i�~}�:�1�t~LYZ�'vq>�Z��P}���¸����t�0~ݶ�"���Bl��[;���Oj�N��kxtB��MV�����p��]������/n8�� �T�qP��x�f�'���}��%!����B�乭�.$�&ק0t��b�8/8*�� ��J�ÈzGϯ6��+��<)12����wL��M�g�Ia���W!�����kd�R�9w	y��;,�l��p��2c�b���)��K�TKS?��>}�]�vG��t�8� �� x�}�k�=����"�D����k����Ϭ�p��g�׍*i�[�U<-(�\b�F��ʷr=��7	z�� �-1@(��Z�D�8��_:|>#W�n*��$Z�fJ&���u���y���[1z�Ql�Þ{gf|bbBds{���9DJ��)�׳A�Gy]ܥ�c�ҭM��SǤ����9-\�����hapz��fҭ*�"M��3�� ���̡��f�pƬ�M��^�!�Һ�L�S��oi�t���3�s�c	�{I���ʃFb�&�a܅��[Q�X�&�3IXD�W�WF�"M�9r��[z�������2A��*)�w�̈́�^h́|",����A�c s�\�9��ˈ�P^lp
R��C�^���@��+Cƾ�����\���	��Hn|�
�?�2���x�9��wP����_��Dﲙ35='���>Sb��`G�C��B^����oSQZ�V�Pp.b
-��`��%�����*����b� ���Mc\5���[12 �S��l+���8kQ�L��mKowCe3��{�؝��y�nt8������0��Q���R�������fl������qse����SF2A�P��GB��A%^���G}��k)�a�U�H'C%�͞��6�L����g���n��=B�������E.�}�L���Z�9� ~�4MƂW�$���|�����,��[�y���Yc�o2�T��1je}Ƚn\�����DZ��4�׏+qzK��|��&w�I���5�\��]w��pL*lƣ�1@���f�o�O������H&+�f�zeQMo�R�AR�U�Zgm*��3�&�ר�)]�Gih@�j�)�u����h����+������Z��FZ٘�>��X���t�OQq�n|���X.�� V$>����NW_<��qE4���7���mI]��8E����fFb1Va0��,N���P���P� U%�����r�c�S������1ML��X���K5IQL��v���5�(sL��d@ް��_�-T�@rFM���v��:l��`��̼�{1�-�pbp�'��5�
�����ےh^��J���x�WO|�d�X��ό����p̷��|���'9
^<5"v,'���&T��%աo����S����A�$fMܺ��1Jb��vfذ�p@��8�%�<�1�8��S�Vl5A��={��r�:Q�ި;;וǘt��}W�$���q�_Nr�ӈ�e������3p��M'���G�-����A���DН����^_����_�+��~p%��-Y9�T: L+���o�{�������$�4L��+ bT?�K����D�K�������Uߩ������Q�1�;tɜX�{)�4֚X$�$w.��a�VDE���K �#fi�7z���F_����>yv�y�Mp�J�nw(Г��^ �����Ǟ%�*�hlՃ�nѬ��ަ"YV�JhM7��rv��Y��O���ߑC%��}���K��Ӈ�t�3X���\w��xh�S�Dꅻ�	x�K�ȗ���A�~O�M���=&r����$����W�f��SS;6�z)�TJ�A�
���5y��j�#��lv$WG	Jހh��җ������⢋�����flL.?'Tn�6���k�0?���9��0� �ӌ�5�-��9���m��-�2��M$(w�B�dK�D����7zyٷ��a7]�A}���?��D��D<@�J=jbg���IS)�Ck3n�:�Y�T��0�����"�X��VJh�ˋ �1yd
$�9�k喲 �M"�� �l��p�G���/�|���ה�<�oh�2��'�:	p����,ȟ��1ߟӖ����YƗ�{kc��͂}�d���4V�j���l���,����N�
���פ���P�1�eb�dO�&K<[<���Q���2�^W��tA�o���D+��tAO5��=���v�+���z�`�3��*Z3�=�e��F�R�������0Cn<�2+�X���4�f��&�	^�p��{k��9��r+"���gi���:����8z`o}�-@̆y�3��*{�'��?	}L��G)�F��3�<�C` �7.⍕�m+%�M~��(/O�v�x�3Sp����`���s(Y�+[x�Pw���{!��=���(�SPϕ�|��;�����7�b�{�R ט��.��3��B��1� ��9�Sl����e{����%�)��S8_@���G;�R;��K$���Jw��P��._���1�e]�+��w�c�,�{�qH��<�fs�*��̇�Zl6y��N�nL4>70������`:�lPge4����G�!�20�}���x߻**9�Vˉ�g�P�t�+أI< &�~���]�~�|Cm����B��j>ޘb�+�<�v�*k�^|V�Ys���w����+�}�\g/��ΐ�D�?�8H��{��\�����x�B�E�_xU)�e<�ؑ6����MKb=�вrV��)�������s����O�U_�mߚ�*�ܫ��Ô�ه��(��}��ͭJ-V��W���*��bw�Y���$&_B�h�f���s�y?���2������a�K�>���f��g�h��w�ޯ:�ӵ?Z;:��(�T����W}�W&��z�3�J�eP�?/���f��of"��������ޡ�+���{�0���ϔ�hO��`	8�Tkj�˞���K[�ب�@���H��Մ�@�������I|={������]U�yYP�"���?�e`��뒋����)�BCt{v-�ð�4��Ӡ$��x�C����-|�G��@�}�
��@Kf���c�VK��%줯e�,f�=x2FUn`lA e���G�(�i �=�Q5������7o`aδ,����P�䤼{�����8�����`/���[݁�%��*�dM������I	�>�\7���P������(�l%ߝ?����&��m��h�TV㌛Ao��䕀7��$!� (��m���]�C����R$x��i&��t\çwo��;zؑn$1^��uX�j0��8�گ�"Ʈ�hy0v)��r]NV|o�����	G��(+(�^l�֬��s��:1!^���U�ꌭ��D�4��F2q<�:��t���W��u'�:e-�mik�RWs'A�E���ꚇ>~�j;����l��JsSv
[��v�Χ���5��	�g�D�.a��#�k�[O�vG)��,�p��K�C���hp9���xW��#W�l���5���@��l�@�����T�K�s%�a�����Ü��.�PK?��Y��1s���ԣ�fY>9^H�d�W37�v�yH>��`�[K����L�i|�L�|j�,���N���� A�
�]��������f.؟��v�%���OS	
x`F�M�2mV�L��U���7U5g�a��<�����C�l��'|�g�S��+{�x9�<#��u�����PHH l�XLPk�vp��T��l�-��k��`M�Ԕ���x�2�@z�o�%4)0�=�����I|�`S�YQڧwkC�
�:DD~{�A!-��	ԥA��<H(
��Ű���1��Zm�\�����}�V�,߫ �����Qej�j[P#z�ӈb�D�:N�q�+L�ȱW���$i�4W�.�QFe��n!С,'m�뿟�O���U/H�c��З�x�Y&HO
��j-�	����>�T�-�Z�2�W�g5��,��b�f�T�;E��7U�GUφ�3h�t���,�@�<����Fladq�BX��GҬ����9̩X@k�g�D�2L��t��b_� ��oj�s�.�l��7���Y���8�H�Гn��"�0����(u3Őe����YJ�;=i��=0�΁��g�-��l��9�Lf�t����V�$�0���S�r����GW3�(�R����ٞ����wh#���l�Z>����$<V�e�[�%rD%zf���X�0��PK��'�Os񸴌��/�d��E������
's�Ĉ����Ɛy�7�l�.6.�sJ���C�b���|�0}l�I�l�ۉ&gE*c���>x@~�� ��Iu'q�ZH�x�w)��<�/_���pPv�E���/0��)���|��/d�*���r��A@����f�*=�=ߘ��p���
�����R���O���O�9lS��g>L��2:�]��q~ޖ�~���v7d7U�G�ɶ������'��&b��g��7aě�zJ�\���=�nKt9_���T
���Õ�X�j�p�o����>/��j��.�O��d��x#��m=e��g@\ ����و��쪫)��Y8O�Dm�ϧ�Y�q�9��`�q2:���_ �<j�G��w��V��<Y��ʳ(ɏǽ� �֎�i��`�yu}R���W��#D����<B�Ph@	`�i��Bg�&����
 "ܱ�Om&�VA>^��������U��+в��G6��0�JA b���y[S��ȟ��:�w�C���bjd��)�xa�"ݧ|��}��ٝ�+�I��g����M�b�]x���5AE������%˰3.6�ٯ�_D���[��o��B,��H���{�q�v޶�c>�x}�ߘ�	�K���;���8z{��J��^ �Ōl�6V.o��8��ң���o��%i{���JM2�PŰ�ۑv3+��C����WJ��{l������q׳����K��	�#�P`ʝ��u�)��݃��7� ��w&����w���^�u5M�a&�S�� � @M��6��Q��P����+|�~[����Ko$�Z�PH�6�,:��*
7.���#n-ۇ�4�=:�_�]���HF��IgE��l�.q�;�Ş�nQб��,<|�k�C�%��*z�2J�cgJꓔ����$���{b!h�b��c�o=�6Q&@���[�Jg�����2�d�����R��M���B��RN
���ϭ>4`�P��i){Cow.�p���F.4�`c�0sʪ�+u}	�� '��������+�)���6�F�A/R�j��fJ�O�������s}?6�I��Nz�'����LNC�1]ŭ�iRb���5ij��!����%;�(A���mf���r�v�`���'�j�F������2Q
(�b=|U�v`	����t+3X����g{/" -��7r�ʕltӰ(;E����������;��F�̖w���1��_-c�NL��=�O����6��;s0<�ԗ;ד�;A�R��i��i�Ҋ��tJa)$Ī�)��g��S#�6��9C/IL�zoF���n�ȫ�A����іz��~�~������LZ���ɗ/>�Z�%+���3V�h����C��%y��eG�U*Y�����x�W��I�l����6oQXT`��,�!@��T
zk���I�Gk����Yxֺ������cLކ���&��&�Î��"9x�3�/�0C�z,HD����IQk~��G����K/zh�0�A�I���J�Pv�Z��nV�R�LҴ8��"�h.�x��~A�¥u����Hܼ���6O�:�Z6�f4J=I����|@1�K���ڋ����<ؠ�+n�	�Lh��g*[��Y���ۦ�F�{�M�	1"#��Om`�nh���Q�/�����c>��<�( o%��0�`�hߴ�T>yj!�(ow�&��TՌ׳E�-$�t!����[��<���=��(3���>�D'�c��li�#u����X��=�Џ���/1��dE�eT�X��Le�B'���4�ӄИh�D�X���΀7&W���j�W7��"�&���|Acj4|��ͯ;?�ڳ����I��x���s����k\�{e����� �
�Fؚ�[�x��S�߭e� {ѕ�4Ɯr��k{%���b�ϧ˕�y�1cL�+��~�����B�FV�.r!�M�4�Y�z['A�N�:)v�#�ŗ��~���2�_[�Fcbb\�z�����,dXPv����C��I����5����L��P��5����k���5Q��Y=�s�&�ԭ겘�ˍk��;D���A��֤���^�rz��1[-U����k�
$>̇o�!�p��ʷ����U���Ͷi�E��A S�c)�Ay��!f>��V��B�ܬF+�R৻��{��u~��7~�$A9;2�z�[�eO =L� ��a�wv�sRa���f�<���T��\�Z���r�i��\�/8#kM�s
�9rЯ�ʹfdȠ
Q�[��P���� ��:�X���X~
,T��^�3hh�90qZ;<�J�- C�y	S�R�Ƀ�ɩ&л�L/I���%1Zб1� ������:j�x@���3�4�����
9�D���)$�#��Ei�����!���a�@�_�[�ۿ��Ǽ4���]W�`��	g)�i�%m6�+�ھԅ(N`�7ʚKU�J]5�Mu�i�R6�(�����eI1c���8p��F�J�����u)���̓ECЪ�0k�Ґ��r����Ω�G�:�%���&
 ~�>�ŝ}ME�oiy`,�5�ozN�&��'GW��l
�ڐ���EU�"����+����j���<���3iX��9�~��NU�	!��Rx���H1��c��f���j�H��\�(04Ѱ�v.Zrrqf!��Z:�u��#��;��.L�
	>G�+M��o�.��au �u V���#!@�i0��s'��s*�i�tS��ܧ���&ݙjj���R#�S`yP.����߿���n��ll���M{�}�?O+:�2�&
�	����5�c���ǣ�1&�����+�MK5������#[�ʝiX,rzl�Ke�M�["��wp7����bB�ei�`H��Hk��9^�F�+Of�{K��?��:��i�ϲ���M%���*#G��`���&�<z�L��Wb�j�xTT=��m1F�[b�9�!M" ���p��SYf���g��ИlF�EtR�3�{�,<s�R-����l���-(��S'�ה�Ip���}��g�3�s6��Sr�������:���<�Eb	���1Ϭ����&:���O"���A�?+@5���L�/���2!��JU$*�IZW�5$r|2�>n�0&T��
0��y�7rog{ݺ#E/�Pa?;��T2^��a ���5�K0?�ql���t;ut'���ow2��p�yo�3� �����Ԝ�����yd���u�u�J>E��,���qA�e��Q��i~��^���ҝSۀ\&�����͉�Ķ^�h|���[��u~�# ;�)���
�'�����!/W���-W����c͑X�n���㏵��Χ�Ŧ9��X��#;�{��/���h/�g�g�P�3������8�G����L*`k���,�������ˮ�9���1�y�ጞ�׵g�����*��
���1�m��Bq�^�l�������ώ���ۅ�w�m��D��6��E��14�2�F,�3���ς|;�F����'�7�m��_�*�#���F3*��2��6�Ӣ�hS��I놆�0BC����x��@{�u�.eh�����嵤�T�Mp�Q[QXd�0�l�;��[U�L���������s��F-���|���Х��\��B��������`����D������6,��*Ab�.�������
�[����`Z�ω�l�ݸ��\&K�tS{��4�V���α N��]���m5O�v��T5�?�!}��8>�-`��&	~��+㬔W/tF�p��9���7'ւ��^)���^���~�����e�����~k�?�w�R�������c�d����Жb�we��X�}R�)��@��a���@������Vs���$z���9�,3Q��	G��*���|ֵ�cR���sb�[-��ر9��s�V�T�D�`#�c*��H�~"}*Cm��#��Տ��w�;��]���i�ш��x[�1�e��r����K9�%��2g�����;�Yah�=�j�E���I6�� ɓ��`+������x��z���/o�E�օ>)�A��~�����yV(���`0��}�;�5�[��uLyv��t�^{�k������p�W�'`ۛ��})��մjm���0�"�2���e;��Q�m�n<���t��tfXH?�SN�����X-�*��f��KE'���
]W�-'G:M��B\�!hP�9�:] 롥 zp>�:����)h���]��F�|ҕS0$�j�]47�E#��g��>z*�J�sk��VQŕ���n�̇k�!:� 3�	�;s�
+�$\�`���s&��H�z�e�w1u�`��Q��˘�S�&���`)sӘ��K��kn�cFDF�vOh^Z�2���)٧i�]�#@�� g�vc%�JHvu�Uzؑ,��R}h:�r�v�on{���p�!�jȁ��*Y�DAy/Yag4B+9�"+Ϟɟ���N_w�նl�!����
"�j�>�3�x8�о��∺/�_�8v��+h,�'�r^_���u��X��{&8�>��y�@�K�������Yf[��X6&�S�~��K�@X��!�jO��N^b�׺�����s��Ĭ�Y��8u�(����تD����I@(���5��.%򎠌V`�Eۋ���:FV8��cY� �k�p#@Ƶ����sh6d)F�	��}�h���^�'u(�������)���^�����^Yah]
52�����
rK������E���[�	�n!o5B�Gƀ�K ��;��2�(�����<KJ�5/�i%�6���U���F,���<ژ ă���9/������Ո&d�d�54qt<��%�q(�Y����.b��H|��
��ęi01�9)�y��n�Js�3I|�K��Q��mͧ6�D5`�[U�~*hG���a�ev�jZ�q��tk�pQjz-<ڃ&�$9���?�L��j+r7�Uv�@�;#�JF�0�0�㒒����n�=����]��js�JC1�%a����PS�l�dz�#%�X
���%��C��՚�hWt`9,�t_�ebzB�j�]�1"n�'�s�,�(�����-l��V�����=N ��9�.t�'����.���o_�L.k��<ȭG����
`v���a���z?b��Žѐ���N��م)���U!��k��s�ˍ�[8-�����o�4K���q;;CJ3�Ho��F��q1��,ڒs���+��_���O��]7x�N����{SR��Jt�9N��$Y�\,o���83�@�+.��(������;�[�aT�-�N�ɩ7��?qL�Gy}���9�/��?|�����'m,͸�_G�%��'7�m�Po������apg?��3;O��3��ܘ����D��4��0��a�����H�7
Y�3�AQ1P���j���,һ4p#�N�����q���q"J�-�n�T5h!��M��{I�[�k�	��w7�a��ڽ��어)���9��0�B���hyZ��6S�o�ĭ;HH��l�p�W}}�X��	.RpW[>�{�b�dTa��aL�w�W���@rl �d���0S�,�LG0� x� c�s�L�'�a[x�-"�$(��J�����jSҢ�_U�XI�l��?��d i�7-٢X���QC}�%�K�9��ˋ�	>���B��"��<GgH��ags		��R��?
�PtTr�ul�sz�V�� ��G�'�sjK���S�o��{�<5�C_R�f&��~�>o7�� �]q�q��Ԭ"u9�2$��T�'�ָ*H�~C��h�E�V�[#ȄU}��Ub�� ���G�S��mi�ˈ��� ��ź �e�>(QT����U8O16�
�O�l���o,ԁ� �8R�}ύ \{�1~��ZY6R�m�t�gS���V'-?��3Kz�4S�A[<?%�#۬���PQ���a6+�2��*���f��z����aH�!�_6��D�L�ԑ?圼r�S?M�x���L�-g��Y��@�S�Q�p�q';J��H��Bn��	���%��E����9���@��2췛t�}�[�]L3�֮.��3��fS_��9c�%����Qi�J���7�Ku&��Ʌ�CA}j�
'C6Ocon#0�2��}���ƙdEc%��:<~���.f�"�O d�eN{��A�����W��l��G��օ{<:����[��W��3���6�U]�CΓe�k_�-�,��%�<�P�8F�0��g��X���՘�)M��뀪�Q��Ah=�Nt�ɩz�u,2t�	~�i.¨�'uZuR����v��\�#�N�UM�H���lF�B*wT�T橄����"�{%�ȭ�����o���>��/0�i�QA��K�1��@�c�9��e�8�'`-6�FiI���dK%�j�\0S��,�WEɌާ)���=���__bwu���^�Laݭ��ctZ��w�bw	0ݹHHqQ�م����i��'_��q�����`�&������VMX*j����1��e�<�L��k� �?`�7�\N�*bD`WM@U��r��ij�9�=�շL#��mo���\>���w����ڝ�D�y��ĴXG�N���L�!�p�ۓIr����S#P�7��^c�T7�niQT3�����
)�9E�W	��:Y��4��f��R\uL�ߦ��b�r�(�ROU
�=�%Ю�~���~�˶�>�j�ΚN�;�8���0�|�z0b��sW���Ϧ/'��'�6�e
n9Jqo�H��Od��8p��ψ�pxV��Ǐz~�7ꩅ�`}d�6�c���ڸy��KT��r�_�J��w3wt�֖G���E2{
R�K58])�l��K%������� �+c�I��y/�j'�{�	�� �T(��[#�`���PT4d��BVC!�6
/�+EI%CZ�̹w3� �L\tE��\B���u���9�l�\՜��!��b��$#�o�}\JC(�?I@?���M��%~6X�_����E*z�V;F�����-S��\�]J��B�<�ѭ�?3����셳���30��	xw7d�G�naڍ��S�Zi�����z̈́A�c|Tj���`3�Ǐ��|@9�]m]�r]�y(7B��g�^n,�:�"��q�iA��{3�J�'�Iݡ�;�pQ��x�u��o�o~�m|{%�6��¬�@0q����D?��������fK8d�g�<��`x��˿��G�����=��@z11㚃�iYqM�	~T�u��Fe�U5��v�֣�<�3��B�yB��AA����͵y�q k��l�����h�!��:� �wQ?ηq�I���ģ�X2�y��ڗ�ϐ�;��;aT�%/���7ӝn|sL+´�S���g�͞؅�터�Y�x��'-�ي2c�W��ǝd�Ӕ���+��@}Z�{�(&��)�N�Z�'��d$92���xu���z#l '�I�R��ў (H[��#����|��Í��t֔�RW"m�6�V�?+O5��]*��K]ސ\��&4���e���G�����C\y|�h��X�Q
]�=��?����mZ�f#:3�d� ���EM�=�s�>�H�p�@��~�M�Vw��hDQe5��B�T���&(�m��d'�����#�D�|Ұ�����j�#�Ŏ!	 b�B�FUfŁ�Q�5pΣqI7$<=�аqn	ߩ��,>�
<U��5��m3�`7(��XO$��@j&�	E����6����E٩B���l�Z���E3���k3kk�J�uő���S7��'B�rX�7}�p�3����b%�G�ц��N�N�:��E��# *6��	�O"���2�%i>�g��o4@Έ��Wɽ�_8�����X����f��:�U9�,x�����+��>���y�Ƕ��LR;��͓*ޒC���F���]�l؆�\&�jA�B1G/�E��f'��9�1K���D-�M�	g�ג���F\K7a=v�Q�(�z?B�ʻ��"(r���v�N�RP�a3B
��y�e�|���R��!`��z�H��H�~J�������z0/A�N�¨�Ŏ�xIN�޿R�
s�|��ź�f���]7^ӄ<-o�#X��}�՗��!*� %p�dk$i���-o�44=O-5���:4�"T �:@Ed��ک���+��x/u�"NjN�<���:��D �յ�,j��t`��9��J7U�KG�*a�΍�+lm=��m��_���?����p��-NR�O��I�ݎ�����Z"��r/�r��;P2�Wnץhw��sb�S�f���7K�b㰇�������=�����9��R�p��,��E�H���|�S=}�,��~K'���i�f�%Z���o�ր�ē9����(���Ua��
�3�K��_
p��n������'~�'����s�7�%n �:�L��b�h�Y+'*1T������:d���&W�n�){졳g�Q�X Ņz�������d=y;��v+��ϑ�5I���U���V�n,Ne�K��������i��P���)�����V�I���T�ď������gC���r[;?��2�k�0E֨�Ĉ�R~�&�T���V��ҟdN��?��ӫ�P�9����!��+T�������c�ΐ�t��s���m#(n�Ƕ<���'B6Y,͉�&���s<��H�]TE45�P�T�$t�����5&��IZ>,����𼻾�k�b%�A����y ��@ь���ꚪZ��a_��[�O��zcL�鏤�<c�\=w�xF����.�Y���&�C�y��o�/�wxn��r��r�@sV�S�2�4���%Bx\,L%��K��M�G�ok��Q��{��W]:S�y����� PN����G�Q�}�y����� �}m�� �6���I1�0��j[ۋn��S�=��e�6���� �v�r��J���U�\���$$�Gҁ���wё˽y1�CX�I�s��n]h/f��f�[�*�S�3c��v|���2%�D�BKJ��%Z?�TPY��J�ғoL�p��G^BkQ{b���X>�>)�LB9�j#&������Zg�:g���f�Du��>�tݽ0�����:�!��C��H��(�����i�.ť��(���j��~<#�2���Ǳ�4ig�0PHdnX�����5�̪Ngvd8���*�wh`>�`kL���e;�	�[)X@��b�ߨ� Az�kd�+�f=�c9�6�*��ȧ{9$*T���,��y�s%(g(ʅG�Z_�ꌘ����A��Wf��f��O4��޻ʳ���ls��%��7ݏM���ϗdH�{����/�P6����/�÷Yϗ=-�)~!?������8K��Ku�c%��;�05���ai�ftB�۷cO�x�Kش�u������a��I!�W��9w�4�-�������}-�H[�ӆ�=6�����#�@��C�
���S�K�`�[`�)�xT��۝5�j��/�0飻�kT���[�x���
Ζ���ɞ��"�86k��a��[�X�e�Gb�l3��Ԣ�+��/~QF�YM�-��i��a�Y�u�IXG�O�s`��(JT6�K�Q�F�Wq��=2��{G��8�D�<��ѥ~�I{��������)ww�Z}�'�n�QJ�AL��V�$����+yD�ʒ����ooy�*ݲT�����_���Z?��8��Tk��w���[�L���O�JJrQ���z�6@�������������)�]����cnl9,b�՞�X�i�L��a��(T���� ��	W�q^�V\?�	�s���7{n%��M�*�W:�h��������Zљ��?h|db�3����ߴ%U�GY<������#�`))����lW������񼮇f�?^�t�VѶ����W�Au��!����U<�ĩkM.l�Q~���ܼ!�P#�A��~lש��x�)�+aci��;QnLv�iF�0.|�SB�(���������\d)ʗT�c|#.�e-�xLπ@ǋF�+m%��{b�����p	@
�^Y��c�y�*�>��ƈ#r���o,������S�5�ɭ��{/�����x-������r�Z]�a�Ӂ#>lT���1��bg�#���?��,f�}����ؠ_��b��ۃ��%[�Mo"=�>iᣅ�e̷�3��M�%�|�0ٲ�=����X��RO��cC!�.�9i|ɔ�ȉṆ|j=��&q?��	n(q�mࣂU��l�s�d!�N�~�ph�ŅO�����M�(�V` _3o祧��s�481T�����k	���)VBψ}e`�7�gw3L�ޥ�V\�0	��֖��v���K.{,As"���R�%}�w�
{�t0(ǳ��ЙUHy7���s1���߫�O��2�|�}�^��I��}����o�}fiW;� ���5�&֮)���$��z�_��{*qg�k�W�*J�fT
t�M��]˙��	��K�����\��8��}�G��x��,TXc�^�Cz?�~er���7�Z
���^�6~�((��pf��^��w�9�r�a�o�;m��<�Ҡo�!F7<�c*SA�M�x2����A_�<m�;Z vi_��}
Fm�>,O��y��� �UFU�;���!1ac!�%�����1��gӠ����W/�JFS�E@ۉ�Gq�[�<E?�y����l�~���ƂC���6��e���������%�oUl*�=��~x������b;�Ɍ�@��*uP�iْ����Z4��E������MpH<OonZ�jdDf3�G�j�!}��)�f_���R��NZ��G9h��t��9�H������U�S5d��q.�q���;��>w�臇R\r��Y�wm��P��Z�K�2���D?�x8�|��$����S��>¾JA� �.g�8���ɀ���ˡ��ɺH��غ.�UfW枈���|D"�s��QӞ_*�C�va�����d摈�B��Db�2Ht��1��.�;n�Y��p̖;��^��8��b�v.
<������=t��T,Y�#?�"�wr|ZWt�k��qMJ��r��Z�P3�i�?�҈�	����X!!{.:�-E8���)h8o�0Tl�K��W@~��A>����ƌ��,*Z�����&�b�=�{u)"Bew��;!>��~��O���PP�(�} *,��/Iyf�8�C����8�m_�>�ޒ��j�Ԩ�\|=N���>�?��?�"*_S(��A4y	�*����MRt/�N�J�����>_�P=���gV��e15ש9�{�;f��L����e�ؙ���؞��T�!�\��=1�)��o�5��q�z�1!���Z�ϟ��%�aF��.v�p8
��>�X��:d�B<R�VGAı�&�����M�x�����i�>��U/��~�1�g%y���U�!~G[
b��9�"5B����*�sɰ,,���NN�s;'���ሷ��y�y�h7�7���>��<b�C)�*Fn~����/ �»�~|2��h��}ؐt�'�ks���2��Uw:�~�}�]p�e�'ĩ�k�f~�%��ӛ���_H_�L[��Cq~�o����#s��HG��������1�,��S2
1�1Z]��ӭ�e��5G�sf�s.���P��J����Z@��$p�!#�i�J�J�H}�X���j�k����Lt��	�u%oj`��ס�A➶lt�V=��*L#�"��.���xT:afI�\{�t�!�U�\����B���|(��ip�"��.$ʬ��v�&d�7��LۛDǹ��Q�	>+x4p��jR��U@b�W����X���մ��MA�b_kQ&���3��爤�h9�E� T��~ѱi;��������ѡ�Y�zt�)e��=�� :,x�f�~u{���� �9m�\���PMx��ZQ�o�m��"��7����=�"m	���?�t�PF0�C^��߭�6T������lc�0�P���E!�ZuC3�M�SڊP��� M;��}���O��>�\��/���G���v�]Ѻp��aym#I(iZEv��i�;|l�	<~�OR[b��?���rFG�������<Ѡ�X������jsP$���&Fp�ȏr$�l��-&؁��u͑��/�9aH�Tb�0���h��t�F> )-� �b�[����*�a�G�VL��9ʶ��V�T^���w;>x�!\I��K�7���F��e�0uv�$(�T�Q��!Xv�ܣg��;�y�&#��@��j�1���;Vt�m��d�X�V�"�����Ӏz�^�!�E�%��Z�U��7�%��=�̂����Mma�����!jj7(SP;zMZQ$������[�IHlݐ0���~��[=��,\�����4oZ��ζ�(�{�Dwt�MHC�+�KX`<)$�]�?����M�WwD��mQ���v���ٍu�QR�L_f�O
���O�B!�X����1�p"f����D"+m�oH~J�p���uflgA�g�`	ɓ�
))�Ϯ��S��wk�lF�EȚ-�j�^
kѼ?�J�Nԓ�ᵩ��yQ���Uc�B0��4�������!J`Őv[�F���]>�z��Ĺ��3�*@?�(7-�bs����eǹ�<�*���||���8��������A3S%�m8I�v����KٗU��զm_��ޘoT���N��A�=� �Q�7�@j�9��$���c��xKӝė`�@�����\@f4�d3J��`2��H���uR�'EG��+� "��XG�R�����G�zf@$*�L[f�]�.��Eo��Z��H����Fm��}b��/�d��J\�I=e�!y�0X�J�g����f�>*���E�9�zG[y��Z�E^��"ꮬaW�Ft����R(� �˫���I��~G-���q[_@DȽ���n��~�c:ƈ�gEժ����d��q��;�w��?��4:G	[�؎����m�v''��)�x3"�/������]OƆ��
�'M����� ]ջ���)��t
���vc�u[����ÿʬ����1u�@V7�	�৆���dՔ_�Ul.."m�tWQ�T>c9{Q�IM��Z�9�h��"�׏�c�	룞6t7���9?SK���h�P>X-���_��A������^�}9�92ͳ��F�h�9[bE��Y�����{�_5�z��t��=^v8V�ӡ~W��{���3X)�t�Ȩ�Z��C����>�I�"����f��J7�=�j+t�'$���S�`���b����N���]�&M�!@N����@��j���/1���T�'�R������ۇ��E g����c���A?v���h�F�����F��ɬ�$��j$�*��NC'e����t��$	�e���p��͜����Ab�V�
�Xȵ�W�N���Z�V�OOrd�3� Sp��%�>ڴȨ�!�=�,��_����;,�µ {��q6\���M���E#ې!.<�4�Ȳ��
�@���,��N��?��ҿ��a����I0D1`��+�;{4� n�9^s:��.���	{�n.��FL����>�B4��J�y_	9n;�9?�#��Ke�)G�� ���@�UV���������V�i4W�F�K�1 �b�a�f��Ӫ�u�gdU]�@^��9ۯk� ��l�T"(*��*sT�x��r��U�����΋�e���#{�v���b��`�@B��ŀ^�~���Q�5;
��bY	=Mk\֕E�b3v|�\J���,I52��@��&[x�3˘i����+�V'v"yw�t$`o�L��g��| !�V ��Z8ݮ�/����	˽Ѫ��{]�W�Օ���q����양��Ph'�Z�r���9y�g���W�Ɛ��ۻ�� ԯ���rv�V���o�R��9I<�(��Q@�����9\�Ūo���ǆ�t|Rσ�2��?n⍺ŉ%D��g������Z�4�5I~�65PʙkWM��k�׼a�O���d�����a�|sw��5^f�;@�'ů`|�bk�Y�\W�/�`�d��Q~�����z�`�!��,Q��՘�{�2�򧗮��;��.e��4������
���i�Gj�bg"H�F����O��AQg�㿘/k_Kc�'�l���So��Z>�Q%2dt����K��Gw,Ț	E)�n�bR��7\�b^����x�a&�d�U57�v���P�����A��>��B}����c׾Ӄ��@�U���5W���g�:��f��Nle��W�Os�"J�P�ד�}�;������{�Z�n�h�%u\��������+�������m���/����@�֠��:���Ȉ�����tR���]Ե.Z���9q6�~��fm�[5V���oCw�������sAd$`�o�Yh%^˗��n*k��c.�=�lL5�?1-�{�+��$k���'�n^�cUm��P�h�q��F��:��y���K�0�<q�^ T�㏖ȣ�R���BOҲ����&�rxH]���5�M/���'!I����i�q�FGR��|��W�r�DnF��o(�9��G�b������.p��ހ�XR��?��U����ҽ�&��y�$�j�Y��t�
�c�ט�|~~�.�O�岑��h�`���&#	�~8��u�p����6���FI��<+C7j�M
EfW���)��S�		s�0Ϋ�v/� ��<�?�+¢�'��e�5��v���c�2��M@I����qI7��P�޸a�p�z��g���}A�O������U���	c�w�@�\<�����Ɵ�b~W# s������e����4�b�H]����!�*:ѓ2�զ�aL-��B��m�ّBI���d�٢�I���$̉�=ց۶ǃ�AZ>��~��+�_�r&��_���9dQ֫�I$��O}"g�9��)������]�#7E/�uS�Ԩh�z��
�L4�$���4P��WqgJ���B�c�dl��d+�җb�������C�-������rP��}�u�u!�`vB ��;oP��\:���w�7h9�=�)��q`��1��}�X��*$k��>o]���ڀ8߬�gn�mA| �
�CB���$��y�.v��f<c:k�
�K������֨E������Պ-�I��*3�R�ņ�! ��2�]g�7l��,�D;T��� ��@�mti��AВ�����E��1d����o��Q~��#8�]}�������4�y���x�>�?��	HO}�^K����kk��_H<D� 4�YJ�q�K����0�����h��3�zWAtJ[���ter9*Ո��$����7 8/�pm�Y���p��j`Ue�{s���5�ce$�k�c��ǘJ�l�)c�.�Nc�O�]/���c�Ӝ�vI�O'o����� ����C|$��0V��U��9T)nQ���[�+��ݾ��x�Gq����I�FX�~ tT�����$�U[Ք67��&�`JQT���Ì�����b�����[#�̬<�t�Yq_ҙJ�� +b@�l}�-g����|;��R�D']!���:YHf�bF��E����o����υp�s�M�.��?��-6屻M풡lզ^���2hĆ���ӆ�:6V���͂ �>�!Ɠ����$L��o�1��x�~c�1`0�zX��~K�g^ѤF�r=�]�1.B����wϩꛉ!�����Y�&Q�
α�GVC'������� k�N���k��&�8��C`�bݱn�z��Ւg̶��FR�
��в~-y2� ���{�T(q{>��M���Hp����d*�F6:��p�����M[N�'�To���j��P+Oz�lÆ�_��8Y�1J�3I�����1G�hv���6Hq�C"wǠ��7�h��#��A�+9�]��[3�K̈́�d�ArA��RC^ml0R�.�+W��C��aX�M_(:@g�=hs��W��I�U�Z�i�����jt_�}�{y~(B<��jB���̀�6N�F�DvV{���׽{�kIy?f��X-[tyu9L�v���9�T	�h^�ę����^���)�wڱ��B-J�ֶ$o��;�@,h8�.΀@�G?:���x�ГR���28��R�{���p���2h*�s��)t��E�S#���p~go�ғ�EFv����M	��P��[���S�ޤs� 6��v�n��+o��)��ť?�n��J�J{��ڦ�A^�h'�����^3J����Λ��ܒ�=�:��`lP�.�ӗ�9d`d"��Lm�\�J���I�BCu:2�g�����4����hS3j¬v�>(�i�-�F���l_��OJ�y��
�
�*5����5X_��)��������L��{��ZP"&Χ�LfR���w��k]��r��s$Z�~�s��è����t-��ho���Z�Hޖ�(Y��Q���jD$= ��7��j��rEwHYa����Ϣ�/��O�E̚iy�qk�X��ѕ�vrnn���+q��'���`�d^��:�_�<z\
p8|no�rc�� ���iZ6�bv�c�ǡ虁3��	ā:��cj>��$v��<	F HY�:�hI8��i��C�����n��5��i`hGzZ��������� ��bE����i���U�)�� =�eH{��k3C?��S})�բ���2'�����U�f�+{;n�Y�� iwpB�o�����]�����O ��\t�#plV�����N^��@)p��h�'��i��j�O=k�^�D<����2�!��"8_6�����8lue�o�4��k�*�*�	�ү4d����`��Xe�ܔ�����1�o�M��?X(-.#����h�"�ǚ�jԪ1��R�ߞKn���X��G��m�Ƥ��T����g�GgF1�ϥaX�D��|�"�s �!���t�|�";�S�8]�1��+ʀv�}!��Z-J������� ���-�4�W���uF$���d�v��@�����B@��g2�\"�Rc�i"�v�����(��g�w,UI���k��
�I�K�Y����-j���5�m;����P,�.q��Q�� �(+W¯��k�ux�'a�n��]��C�w�^=�XMJ�$�����B!����2���#}���H�x��z�Z��i�G��	9�Rޭ� �ƍ|S��]�������*Q"���gFw��k5*O���a��ne
��q]af�s�!E�"������gJx(��X�(����XK��`�W�m��?kx�����z���x\��7�e2���TS<h@��1�4�r+.G��å�ݪ|���zo�UR�4�� @R���R���z �Jw�Q/�G-<��9 J��Vt꿻f�a�+�Txc��������j�[ʡ�X���:�*����MN�Lx����H4�C$�����w��VXB`ө����|�ĕ
^_�&JM�ī�"2�\ؤ��ɰ��n��agd{99D�&*�'�V�U�9�e�}�?bI+�ٳ$٘(��c�3M~9@+^P}ܥ�Ϋ2�H�g���U=���RJ�Z3%�5�!!ݡI�)4?�"�{!��d���ĉ*�S0�A\N�]u���] ݌򰃏zn�>Cy/;7N�X�Y'�� �qp���@g�v=+�b�� FHJa�W��I� Zn(�|�D }�[��5�����)�h5�1�u��� a�3����J�P6�{����<={��y���%�l���忋IL�xB"�V`��P��h���<��L������PR�\n��,����ɑ=��M�k�mmQ�B~O�ަ_ؙ.�����Z$Rt�#X�T�u����g�~M��Y���+യ@(��w�i�}��y�Xȁ�u���,�ǲ)�0�EJ�)[c�W��������y�<b�(���O�l�����{���g��C��[G
��n�=�^շ3���}\���G�(��@�t&�U&��<�m}�v��yA�ҶS����8%����)N�8J%��z�p1PA��S!�$U�If$��hD9E��ڥ�F�ㅼltU�@�a�:��{E1iq�� ǖ�:�
K>�ݣa�~m��6�`�7)���Y�bM�Qcs��G����z�֝\%�Ã��vF�c�A[���Y���xWu}����E�7кԡkT�ȣ�|z�.�$�~n�`dXzPؿI#R��n1>��%Mo+B3��]��aU�uV��T)"��;˖�R��N S�`xN�yU�@)�t���Ɲ�_�U�s_Z�-ubM��h_XBJ��5N��p�1�Eɺ,X�kd��E�@�N�[��3�����6�l�E���T`-Du �F��u�o�-��z���	���-��~<����#(��
�I:K1�p2���Fju '��;��B����d��] �F�v�y�;J�ք��ȃ���֨Ѫ�qh�&����7?*�՜���|Q��)76"�e�u��A[nz	�h*�����"ގl��s֭���%/%�]�5C�`�����p�BG�q��V-u��/{�U�*�nb�Sd'=0�&��銝e۴U��/����ﺲ�l8~��%db�#j��e�|����);����IH]!�ǲ�ϐ�ݵ��䯶����soY^b7���Pj�uڃ�]�I�mWa=kܕ��%�U��27h�SP[�v�
��H]Y����@k�O�,��I��� /��{��ʤ�.��ޥKE��(N BB�^��
E�og�p�C:J!^�e.�MdP"��p�k�{��@�*�C��A��:
0ST_Ќ@��fd��׵e�Gm��Hiu3��n�ֶQ-��ȟd��t��3�U��2��|�_S��Ka{���R9�M^/8�s��$����4�v��O¡�5'�%L�a_�|������a�[�r���e��Va�C6�Y*���@��}�޺���}�ֳu������6
�z��s/���$|m�&B�b��v��
70��j�;��כW�ӍY6w�)Lކ��MU3¸�=���>*\�����t��\Ry����l��v�O�̤34��=��D=�e���K����J$ӕz�'������-�b��pl)\�%=�I/}H�aa�O8�pu� �qpG)�۲�tb��E�n5�@�̄�_�խC�yUBQ�n��I���9�~�e9�/ ����!�6T�%3��u�>͡S�z�?��9����1v;�����s���,M��zM�&�>B)�º���߁6CSWm^|��P�D6��W�����C²�!1}ۋ~<t���w��x}�E����=���N�# 9�J�j�NPg������H[�vi�]H&���\Ki��)�I<jכ ��kfȸ��_���ؘ��gk/^3��nv��H���|�o�b��qyR�˃g��8��^�*6�i+�  ���(`�Ҁ��;���#��2�b<�E���#%��6���:_�ŋ첚gQ2#���q�f(�
	��;�6�r�?�^����_v���p����e�.�b/���	^���ؼ��8zֽ�����\�ibll۞�Ã ��>=Ռ��Nx?����h֏���{>���:�}�V�dPwܐ�"󪅁w���f�� �o���I����U
���.Ɛ����JTzM� 7,�����z���;N?q}�cC����rXA
���CՏ$���h}��d�_�mI#�j��4�t�]��5pCϓ��߱��
YË�IY��&b�rB-��b�T��O��1�*1��b��[ �U�2�m����$���-�&��I�%g����A�hL#�9��r
�mx�O{ɲ}8����UK����2*��)�+�T���F��!��4M�6hx$y����ͤ���W�!�0�GV�����8�9��h�Eܥ����	�o,'��(�@��P�c�����	�Sn*�N
��$�5���/���at��}����  ���xR�~r��F7�VG���.zm�K	~T]�����#���i{O��X8���s�]�#~��l˽���<��.ԑ0W=�;�b�Z�u�TW�f���<]��j@�C�n��C)���]T+�V��*^��~���o�DS�<��y��u/A�l�Y9i�ٮ��}���M���-zg[��k{0&-��k1;��1�䓀q���gq��R���Ҽ<��7X�����2k%�������,3�|�|}q%k�c�8�G��
�� ��:
�vǷ�v��ƪ${�sO�)�Q�U	���Vξ4�[���:���7&w%ޞ
v�&���e�,NY|��t��3����#���C�TХˑ�H��Mc�-��Y�l��c%���3����v��Mw�r����PPRC����$U�+J�f�sU>����UC��x-�c�`#/S*f���\�I|�Yp�@�_���f����J̏���]��P��.��]�-Ǎ��3}�xU��-�,v��Y��{ ����U���Lg�'f7~��^��(�pU�l�f�Ǯ]�+�4*���f�����~�hp��zͧ�R�#0o�n�f���m�Gٿ}l���-*�	���B���Ә�h��ge(��!C��~�m��%���h�շ�|e�p�� i
`4�_>�"Q��!��t��Ϙ���^�����%5b��ܧ�B���%�}ѝ�c��x�)��#���L�ɉ/𗫤\:'����C��T&tK�k��r��o�����U��n��������&�Ʋ��5�{i���Iŷ���+E�3��8g���hl"��~��쬤�����̜�%��)�*?w|�Ռ�0��i��KXK���j{I��ij��&���$��Kb�30�S.t�������fw-�W�����\mfhPG2�ĠG W�y��<����F}��
�k@�	�9Ne�s��CV�-a�ϸ�@D��W��Ͽ��R^+軱9��V@�}\��zЏ���h��+b�W��4�bѴGT�C�
-��qg���m+�Ң�j�^�;zg��}�\��Ax��S� �{�o��+ہ�;{��?����!������2;�˷����~Q�+V�y'j׽bzK0,�:b�2�Q
��N6� yF0~��[��M'�̗�c��)�:4c�x�˖E�}\9�fȉS)�uE���o�=�:Գ�{��AX�7h~v�׉�$�t���_ �U*�D����nt��.�Z���d>�c>�q}��_-�XN�;7�Z��n�!kDb�?�e-7r�����*|F��`_ۭd5L�B��'�~h��uz;bg���.��/	Lfj��;�'U礡�)=���,'�������M���YF����y�< ���G���bz\,���O�y�?��S8o��?��@�J��"��M��\C�.EY1�J��:3텻b+6krp&�5����ڏ�(�ُ�c}A	���~���Ґ
�g-ڗ����	}YIF@N���Ӗ�>���� .i�D����k}((�;Uz*F���Z�JQ]�ݻUgt�^��,P���Y�f]�YҤ��{,�I�ST�^@�<<.|UB�5�'7 E��O��$4�Da9����[�.
ȅ��^o�y��R����(RZ6�I�X�U�$�c)���QJшFC�_a�2B9���jא3�%pw[�E�>���`J�:`�Q������!&\Mտ�o A�Ad1�x��2�
b����{rb(!���sGD�2������yt�����9,�L]|!��!��A� #���B-i����p�_r���9�n>w�Z�fpZ�&���q2��V���m�~��<B�������u�;ޫP� =(���)��y���8�(�X�B�vT��5��tʌw���`o�Q����]��i]�?M�PlW(�"��b��B2�����&�>R��Mb��β���2���ۛ���j��ڒ����W�M�����>g�}
�Du��ѡJ3[w)OQ��_�˻X�X�����{"g\��|��}ΊVb]g���4���.	Bz�Ʌzŀ/���?��K|X�����8�b_�e�޶r�!��no5ZT�dtT���3�
������ȃ�+8�	�`;r��Q����s�Љ�+d�jk�Ё���P�M�]��-�5T�9u���~�(Z��tЏN�]��{�f:�>Q��z��F��d�ky3�1	ӷ[(-`�C����@1qR���(<�.J⼈&�}��H`�`�'�1�.��)I���7��25�؊�G�V9� V� �Ⱦ�(��ѷDj�$^3�m ��Q���!Oώ��Z9��%�ٳz�)gq�N����Q�>u,��F'(Ją-k���v�C�vEV_��m�O����/\�٢�T�:]F�l��,A�-o�~v��T�U7�|�\{�7�qU&�K�-�q�@�-
��$������_����)���.��{52d4�]ϔ$i�z�ɘ�R©a&��c:�g{��fO�?ƺf�kKU<�+�8�`����#"�kN���Nt�ߤG,Z�JiD^�==�Ɛ�43(�86���QEz��	>����Q�_Y��f�(����Sܦm��״�i'T#��0��_��p�O��c7g�9&�]G�C����-��Vy�_RM��8���b�ϑ:�#�U��k]3�,5c�I���ܴf�����S�Aѯv������#����]��۹3�{]���u��T�~��}�K�ajI��(�OE1�(u�zؙO/��5�*���v@���օ=��	�C&9HM��"z[�}�[_���\ɳ��P�r��I@pk���y�:+��6�/�`��Za�����̼�.8q��j��j�ɑ k���,��b^��|�����g;��
�����h���%@�'�k�nm۰�/L(v�2w�Ww�e���݅H%f�8�-&O�5��Mί����#4��<|�N���;�3l�.9SS�?X�1����k��7��
�#����-�`o���Ƴ�ÒW=ry�u3z��7n���+"cgr�z��|.�r�]>�d��$�G*%������C��i��X�z�l�J/�p�1=C��?�\���҆�PP�G�@�B���O�jKw��Y�b�*�����\�'����#g&���S4�~orwTY7 �<Z6���"�&�(��,M�V5�����J&��6 ���pL|bġ3�Q���R�R�WpV�<.��vwM��� ���l���;�v3
��s������	�)�WU�( D��O�f%�n���Wn�&��|����>�|	��������lL,^Pw�t� J�:�)�Xc��93��I��U���n�G\��|�uo��ω�C�wGx`T\�e�i�D����o�G�=*e�2���h�]#�B�22�'A���m0Nϯ�E�����S��Q�:��%M@�Cr��Y;E��.�9��.�Q�¢2>sp9��м���������4ul�Qe�ѽ�j}�>�uUױ�q�B\���P�n��� Ȭ���۰�����n��`����~Ԇz*�n�}��k/�x-���D7V�y��S�?b*(I������J;>�ọFk�ǽ7���OЁ	/`mQ�B�ւ����Q7�o5,�MԬ�[��ݥ����]�����̴Jz��!���x�u-�4J)�Ra�yb�O�`u�^p�(<�ߡ�N�wڸ��u���.S������O_#gT�|u�� �����{�s�B�oy�h0$����f�բ!��v�P��M�u��<2��+
�jkr�bݫ���'5m[�+F�|�y~�	�U�C;��� ��TwI�R=��7��x�C�[�'j�����p:/D�����l��3
(���<Hw,W�m(H/� G�8�iR�/���*�#a�QH�^��!�j[LN����÷��e�j�pB.�b]=[<�0!���(b�L�f�J�x|u���WUNT�\�b#D�#�xuEcso�$�u0�V��e6$�	<x�rCȤҮ74ة������i��>F�o��y�	r���-��c�>���:$L;h�!/���RfϜ�W��v�<�} �9�@D>�l��gA��7�p#:�/���3��9P@�Ξ�y�[	&FS���Afl�p��n�gJ�vשu�F�o3(5��d �ޫ��t<�0J>�$�`g�ğ�!ch�^��S�UɾUB��c��/�P�$~��%~y	�rd$FW�:[cE����ZH�d��g,�;C�x�_;%�AT G������NJ@p��J���&��>ZM��r�~��^��H�1����}��h��[����:�[բ���޲���7�`e���/~<�бaÃ��(N�d2��a2�0+p@��1��+e��_s�|����R\r����,�}�1Vb�5U���xdM��}��(v��0�
��Xw�@R�4����{��|�G
Y����!��Ty�$�x$�
j\'�	V����ߌ�K���Z�U�#_���mSm��z4�sX�'������9�Bp��ʓ�gH�YpR�u<=�4\sae��G5��� o�q�B�|\ϑ)?\M�����q���F��L"��N��Q���˾~W�R������݈�f��ȥW��+ }��$��,o�P�H�Y�`��)��4q�����)g.d���I��P�k=~W�nAz(	/��10�x�x�P�u\��hy	����p���a�d������q�
��*���ο���/ƭV�h����hs҈��D��7�1�����ȃ���[�#��v���َD����a-$@o�&���zY��F�N8����/X��}�JJB�Y�t����ї���v��e}�]H�x?=_���ȫ+�WA_��j�C��b�0���0�8�U�x�л}��PO�3���y��H�f�(�����S��_ѭ�QSͣ�k������Z���������T�� ����r��B��o�U��1�JI���9���� ߝaD�U�q)UC����b�.rʙ�3<kM:���q�8�>����m[�
11{�g^�g�/�I C��`f���8}E[y?	k��O,�v>�$P���)��1c~(�	�Lws>͕oGqR�L�7]������:�>Eޜ�G�x�w��~M�l�9�A3M��F�[���5�ϻ��5p�]T=<U�m���w�㤁�zAV���5#{�:T��2Ll��G�ƻ�NJe�r��C�tkd�W��J��= �J*�N��Di���m[��ew�P�><Ҷr[����StV�14%�*�7L?��	�x3W�4k���%�&g���:;�au})���/ʋd�	-�A��W�ق�8F���sԜmα@K����nj�3�V�_�"��e[�� �I�|�,��q�Ζ��ȱ��2k �j[�X���ד��d�yA�NW�G*�ާO�@�����,��L��U�۪��&��E&�tДRDe�tCѝ��e=f�� ���A�_�Ook�l�o�̋��QR>p8��.��<��)�T�6	C ��{h7s����(ķ	�8DE����:����+�����"ŏT��=h���)j��r�D9+�*���`<6K]")�Du�"g�h.uu#<��ךd�T����� �j��k��\�V�Y�����~\ra�m,���M�_�*8Hq�6q�c�����N�f�jI��-w�{jmPy��2f�5��Hp�̔!�����HЁ*V��74td�H#��+S�����0��p|���רk�y����C���ف8��t&���yL�nŲ;6�P������/I�E�l��������y/6m�V�~��3�s������>�v�H�=f�������I��>�����0�����u"�w�aS��*�u= ����ܔX��g�y��r^�5~=[+��Y;�r:��Y�}!W� <�E��v��(2t�/��@���#���W{v�o���зV/8n���"�X.c�h��165�g̴�`t>���!(e��{��} �E�������1�����=�w銐+mו�w�d�m�����ck�V:��=B�����Z��"�P�#W�v�D~G&��>�8nU��"Ň�2䄇'�4�/��@㈚ �kn�H8���>X���$R�r��HW���E޾���d<���7O]ܧ�F��,b@�q���~�c|�8�K���.�WI�K�Kcy�E,��`�?_[�7v��~�2��Y��ML��3�\}�!��Z9�Gj�4���k ��C��~������Vp�NG�o�vG���zn�K��pMˍRQ��N�2b�I3D���C����C����i�N�2���!�G5�1��Db�^���j�~��XO�y�5r�|���Հ��˼K�?�d�3���.������u$��7[�b�m�`�k9�C!&����Y�"�%>���v�`~V��QK��L"���M���y�/������&Q���L��ۛ+Ȋa��nC:q���? O��a�0ݺh� ����q���p��pmn���AO2]���&�� w�p5���.���!]�o���l����"���D}jφ�#�c�<�B����B'1h�Ī���>�D���B�=��&�qb���!j�����$B�ee���#�h�(j��벞�7����̕����1���F(�
b���dv�`Q/Y焈m���Ǳ���t�/:����*����ű�m!,%�(��-����xO9���;o�ioQ���۹��}��^�hJ"AGl=�pA���##,�
U46b�r�{0/8�p���cW3�sg�:_-�
��8�e�/=ڊN�:�sJc�HS���ho(-`����D���Ǆ���<�UD��N9b�,s/uF�5�,Ğ�	�����������k�YbJ	*)����w!uRb�Ʃ,�z%�}�Gfa�>��Y�R 125"��0�s�u���S[��T�T�S=p����z�tT�+�~rϢMxh�E|�d��S�o�`!���RK}��`H��#=�+��UB�T%{��B�$d
�ʰ�ebýW��H����V�(ְzE�ȼ�J���F�S�lH�|���Fk�4�=4�j�o#x,[���C�y؇�zK��A��	��H�l?����*D���Q��:�J9G����Y����|'r
�Ȼ6������V�5�e�9m/]ՙr'ݹ����]J-��{���E��E����Wwo5�W�r=���j�Gl�(� ���p��M_�"�d�OB����("�=��U�18'���DJ�&4k�㍍�%z�$�uZ=j8B�0bMx!�Mԉ!8 �J���Hiϼ�x��Aq�`�@j<ܱ���@N4���d��ޞ$35��/�Qh�p��+v��F�:O���e�zlީ���9���
Ĝ�&==��rp��������x 2G�K}U��'�$�[G�GP�@��ļ]Ѭ�6ʸ�p��0�Vr)I~�f�J��N�PQ��V��<f����� k�#�z7�EǱ��K�C"�X���U��[�aFkǾ��>E������HH��QƉ����7���6p�L�ܘ�13H��	�3O�,�Z������)�|uNC1��������F����难�ߐK�16�gˑ�!b/>@��Oˌy�_~�Lr���&�3�6Ň>�%���������Oۜ���2IӨ��V��2��ۢ��s�g}��yX��s���ŭ9t�}��F ��a����Y��������V�(�Ԉ������!�?����(V�n�F�0$��ƛ�)\�b�N�.��7���l���,]7⳾؛�B���opp�ψR��+[��K�>�!�<�1��D�9f��53vhYI����<�)1��H!�m��VϢ��h̸~�WR��b�� �I3Fs�.q�����՛O�X3��A�
vyLH�D@����ld֨7���!e	5YhH�>�86|���?�b�K#�����t�?�$��Ԙ�H�f�B�N�qljĩ�[���c��bRa���g/�2����uNJ�1b��w?����e�UB��V'�$���u`����Obm2��A�\%�t��̽�<e��Z�P�,��P����=6�2�u�������k����r-�f���(���Pld���K ���d�`G~_��at(Z�:wH�2CB�*[{�G!x[zj��
�J�)���G�4��<튎m��<��5�i�������޳�Ô�P������9u����+lZHJ9F��L��k{�o�ת�;�Kp�Mx(bg�̓U${�|Ep.&<kr;��]�r�Q{�U�����>m��ȯ��Y��ů0�Gm�;`3�ZN�
L��arrG�v[%SA([�{��giL	>�[��v[��?�?�Hn2��K7�Y�͎��:^}�C>�2
]�P�V骄a�oY���P����|;�3մ��+�ѷ����Z�����;dt��Ո��>�;[��q��0�LOJK��vp��Yd_.
�cjw�@�h9e�������:��s�GWKy\SB�c bv�-f����C-q�{]�[�/k��IL�$����F��x_��	'ң%/Ҭ+�����b}�̜�S�K.�uhf�����0�k�8#E�烾*E '�i���$�F�$�I���z��iP��T]��k�/�B�b�'���/+iŽ�с��mҧ}%����<���kx�����;�S7@��l���j��B��e�iO1�t�ʠHS���SdM��*M�LVV Zr*n0�4�f�I�f�D2\�u��y�6~����~��Bρ'�r��1̞e�es�8��g�1��Ԯ�/�5V|�.�	!�Ii��J
L�������z�d5�i�kK)O��xL�Vb��l�T��Mx
X'��c���8���k����a��05}\:���P;��a�߽Ï�X߇˂��5?Ή�Jg���	���Li{ ����)1K1�z�Ϭmb1;7�+���C���`�
d8����47C1��$�F�A��"':�+�,�=I�������
�tfftMgQ�����'_r�lpT�GF�J(~xÓiv���:/�?�tl
�}#�����%�	ݓ�����MM��QVջ�w�OCỦ��F��?z"���3�v�/�~~�+їw��07~�1��H��G{�Ε�q>�F-���{�K�n�����
,�]z7]{E�����l]�
�Kn^�;�!'�J�������w�<"?_�=�ȧӞu��f��s~���	�+ �����^u]k���Dv���k��|%O�z�c�r���*�2�s�g3��J��t�U*��������6��1!w�}3_�����qgNۑ�����$ I�4�#>�����5����Stm��&9�E�J+��v�L�9������,�J3.�Mh9���ޝϋ��`2���^���l@�E�_\�?h� ���AS�w�>m��E��I�hOڠÃx���+T�^s;D�at����
�-�ٲ/�&�(HC�����	�l�sꚰFSP|ip�pD�׆ob%>�7t+�'�����i�)�tem( &%���$��G"~Xi���}k@6� �*�Dwў���P ���X&�nL7�Q�QF��:o*�e�($�>��D��� �x�ήwd<&li�ؔ�5��"z�! ��yd��C�`��8u2�.^���^�ɯW^Oa���Q�Nn<
����r����iw�ɲ��=(��˶.1��1j��=��Q|����B<�H��I����s3Fy�W5��YXHњ횽9%��z�{�4` �&�WK���6�v�_O^����5��Ga�R�:���+��^�����_�0U�R��#���0�ʿ#*qp���x���j*X�>0��K�z`��UD�O�N��H��=�A�,Q�W��R�����v��	�}��y涃�S�jA_��Wu��1��}��s�Ja��,w�|%�t��o��0�M�4e���c�푳ÓwC������!�>�d��1/���L
ٕ"�#�H=V�>���n�j� ����q|������3	�:_�{��e
/�7�xZY6�ٻ$L����4r.5kyR�������^�6E�v�\��VP�Ι/��w�����\ "���Vϻ�q���3R|uxX��h���@��ő󡰰+p�
@<�6��U�P���;/�J_�-�B�W؄4���G+m�6�E߲S��׾�G]�|�/�]fSOKf=0
���&��a	�36���o��A_��a_^<��"鞥{�G��EU먶!���5Í�N�� �e���:����3��A����2�mb�.�s��קW}�͘s�ҩz�;�ˏ�v�M�5��	�%w8������e`�a	_��k�tz]�$�gBv�o�?�K+�'�����;i�OQ2.��Xx7Z���埇���l�#t߬v����z��V���g��s�9�Y8��C]�l�;
�9Bm뎅\�B�F c3����s���r��(��Y�$dP�?�ף�	ꥰ#��|ʨG �u2����SoG͙�����p�ɵ��~$��B�"�d_eF���9˹��z����_�����+hH���W��([�;�����e�.ټ8f��~L�\�X7�g�N?��tY �|^��-���ǣ�%Gⲧ�oj�h�W��E�%S$-�b����ךT����[,5���s�&X�}��+����˳�WU��F8��ր�qe�S�Z
a�	�ۚ˙b:	���:�i������H���k2İ�Y����C�ϡ��7BT��b=��N�w���&p�)�82y�,m]-[��D~��}*ȩL�CwJ�qvX��t���}2e�?8��z�ET�Jp��8 N��0��z�?�����u&C=,LN:���V�#U�I n�0��_��>�V��i�  <O��ģ?;�Y\�u7�2�(=��۹����x�e�`�_���0��{���T2l܌#'s�-�j�zt�
�?��;�tA*��
���YYy�g���}�yP�\���6`椱^�YK�GҢ#�x{����Wec|���_eL��~�tLDTfp5c���2�6�dHJ���$�V2�_E5��x��A�?�q�R ��w,yR���o��ɩ����W���rs�GK蚳�`���T�:��:e@���Թ���(%=����5�m+�WJ���%�SA�B<��xMI˥�ʅ �#��]�H������G��.rz���z�����ˈ�K6fs8p(��(�=r�������3�1ct�N_��a�0P��0�����{#a-Q<
�Ը�<�n50:MAo��`����W�[L9���@���͊�:�!�X~<_�zc�(� �r2!w�|��=_�h��%��d��X(/Z�mx
J��&�������
�6�^�u�R}���f��;Ȏߓ����ϒ���_�X�
�N��<��C�Jn8	ʾ3��?^�n�2��Z��-�[2�Y�:��=���|�Tg%$�B8hX�t��-�CXC���_�Q���X���8��t���xz1��Y�G���~A[O���_�k�}��u�e�?95H�e�ȥ�RIw BA����^�~�m$��΀�ZUFTNݕ�[Ϧ��mn�vЙ��G4�6��*�O�x%�/�/�ϊ��݄��kűk T����J��KF���j�?���Է��m Y�b��E�;A����+�Mt�!=i~%��91��7x���io�7��tP��-u��Q��Z���O�9'[1č_]p3>�X�6����3��R�3*�����;[�_z&�@� 2�2>Tf��Ӱ�-Hq� �.��a��j^փ�s��6b�BF�N�9�"����WJj��b6����It��hg��N+�y5	�@,h��d��#���T�O�t<����d�iX���P�0�^��dv,��^��0�0��Lt��yƵr��=e�[W��.�-�j��+Djb��z�i��L��<�Y� ��y�q2q���՛��/���&���[�W��5Gm��Qɏؾ���pmƊL�Ѥs�&�oSC
:z��1E�f��rϱv;���Z/g�H�E�pn�Nnw��g��nT����=��1�S�KyA�auw��@;pRq�� �c�o��q]i����s
hEw�F.�5���K��~�x����Fl�(�۬�'*�D:�)�˿oD��}��7�Yƪ}K��䞨��������%RìA�غ��f����`�I4Z}��?��b*�3�,u�ZǶ��F��I��:N%7mM�-���&��
�����L���;`=�q+ v9��0�wʇ��&ƌ������	���-�1�C���"����ֆ�Ch-%&���a�;j���R�ǂ�5rC�c=��0���sW+�J6��tL��i���!���� 
�I�v9↲��eX���2��j޾K��5uv�$�J���BQp���F��[U<�#?Wջ
�1�pr�>1��'a��p����1)��$�����ZO��������ۓ�N`,�C��&Dʫ��z��W��g@9-f���e|K▪I������9+-z/�FT�U��3+Te��}��/�kX�\����Jf(���[���6W��5�h����v�6����p��ً�W+�������ɾ2����Z�Au�]RSY�Z|�g,|�\�痫B(�ĕ���s�
�:�)���}nݐp�Sώ���&}�Z�;�^���lR(��H�8mb3�3<�A�ޛy�r"�ǽ�!�_Ͳ�J���i;�&.���t�p�7n6�F���,\�Z;���������v�gд�gX�o���S/��_�6�#��[kF���t���+wI/&�x���v?��1��	_�{��1=}l�)o�&w|�������t82$;���7�����1`��nQ�*Xsvy�}��/�ېK
��2��f�:mmRdQ�g���j6�cd��A�Ǖ� P�����ML����r1�o� �<����m� o���^�,�g��Y[?�H���@��8���ֱ�����"f�N������,�d�ǁ�}��K��N�S�t��	<��ZK��HZ6�������lz�9��x��P`2x*��Z3o^g_m�u �ѺO����!ۢݩ�B�A�OLM.��٤�W'Z���O�H�^wF��ї�惦�L�_� ��3�&��W���������/��)`|w�\��[WV�8�Snz�F�.�)���~r����i~��z��_�L3(0��ꤧh��gX�����;f�󅨷�u<MK���j�d��(��	D'���4<Oإ[	�g��8T�I�
t����r���t��[Bg�u��BQ�޷�xq�7��`�gp������N�k��-q-*ee=.�?ya���ϱ7ނ�Q(�r�o(�o�_�@�f1c��˅����Sv������8R[��&���VS��L���w��ߋ�`��O�*��-"����j4q.P�Q����3�����oy�ھt�S��E��sI&J�.�@�<2R�4�� m9�u�]�����M!�W	1M��ߓ���Q���.��'���U�$t�26F��r%rEq�<�"!S-���¹<�8#�T�L�fɠ�8m(��Ő{�	�:��G3G~�MY�Q ���Č��C\��hߘ��!��O�]G0������].@b3iQ@�c�r*u9;�ۥ�����l|���fT�J�R\�Ȏ�է`|';elndu�I���,=-��M:�H��e����[�ږ$<?�l���\=f��L:�ͮ ��3��l��a��LG����e ��CH��*h�M{
�e��!�D�%��`�\�����O̵��ۆo^		� P��xQ_D,8p���> ǘ^jV��yX�U=8��ȝ��d���9
�U��הd��{�W�m�1��)n�4�Lh�^�}��qb	:���vI/:��&��?��Je��`+΋޷�˚e��yCQ�tDD<ɹH*daH0��v�������Ť��"4�4L�A�o��hXw�6ދ���4-ڼ���ʂ)�HhOM��$�A�w���|�-vVz���iЌ�����>���]��i����r�H��qd�8�����-q���jq��� ������y"%&
U�M�Z�y�w��P
�	�C��H�8eN���1�g��R��( ��_��ۈ�E��ޠ ���T�4�2���ζ��m�l�Q��x`�+*�v�tb�/}�2��z$�nlBe}���kXD0Et��X�fq�y�b`ekrG�5���		���ñ?Э>ȈF�J��Ҿ���w��'�]S&�*�A�X<�u6�ᄨ����ͫS�m�q�m�6=dd��1r���nF��q���sYu�s^��17���-��\��rӖA[FP�I��#��v:������bZr����gt6��vǴߙ$!F�}���"��*��b����R�$P ��x��&�K�fT6Ԍ�Ì��H��c��"y��(
@�yƼJۊ�3�\���� P	� ���{ݻ]���3<&�F��_�H���
���"�I;�g������դ������kw�,����F�h��.`DL�3 Jk�Q�P�����{�ib'o-���\z�1{ ����//�qC���[�J���Ԥ��	nX+��%��w�z3fb-߂����U\��lE��j�Vm��x�:�OI������V�՛��H�J�_�)׸gHxp��̃m*l�ßη�r�x=��9�>�^3>���N��9i�ꨚ;Ȯ�� ��9���fM�6U��y���
N�,�!���
�gu��'��ߩ���S�{���dHe���6�^�Rl4�����$YM��O9RPs��*�����u A/�.�R1M��.?��R�MJmx^5r��4���9�R3��6�P�ѹg�Z��s�t��w<��)0��\=�(��MDJ8<C֯�����
6����T�Q۪��xP+�{(��̨�X�ma���ٍ`�"�2�����[)��G�����MB:S$�(�B&a*J����:�1٭���Yu���A&���3�m���(O��ӽ�_��r1E ��%�y�d��ir��j�n	HwDQF�6�1P�o�ӗ�0j���2y�(U��*Dͧ����6OL1�����ܽ��E%O�;o���M�n�X�yͤaN�l}:�%ħm
�s�a4.Ec�\�����27$qk5�wȶW�cG&�U��}x��t.șl�q[h0pB��i�eϋ���8��O��'�co����S�-��֛�+$q�
�8���	�z3����U���W�;/2"9bV��S��Iͮ��J�)Wҳ�QH��S�`M��67�3���=JÙ��#��zL� M��g��$ـ�j���"�4����b��;�!Ζ�`k4�E����cO�w@��<B�6�[1�����p�q��"v�h�`�w�֕��`_��롶�T��X�wѱ
T\q�O}>��i��֥�8i�E�p%oT�~{���NW�I4Ը4�9$��Iځ�P[�&��ҷGڈ)�t�����:x�^h��o���s�"E�7gJ�X��2ʊ�j��D��B�v����#�����Bb������ױ�da^^�@ʊ������_o��r(Aɶ��beOFE���-.���<�����{�+Y���PS�{�Οr?Ęk0ݹ���#B&~�d����7�
���;^N�r)��02Ώ]�ܥ��n�sp/�b�[t��3 �+K��`�����=�B�� �ͨ�&UÕ&��QE���$�l
uN6wO�$�
�24�C��5�QQU�'��w�'y�x�w����E��&=#�A	T9Imfj+s{ꇔ,	��1�B��e�H�!�0y[ �K��nNh���jM��H~�4`��u\z��vL
5='��ۍ(�>͎~օM���!���������N$a���&&(��4�wk���Sr<Wae��}�_��/Q<�*B�_!*tC:װ|�K-�~p��D1�	�Y�h�ŀ���^�CXXc��������bA�^��,��6
<�Z.C����"߹�;��J[��.C	㸆~���۶/�p��֨��a�u���t �1耤 ,y�C!NErΕlC�Լ��fR��y��-���p���=���oU�Pj>�P�Z�+�.[�ѻ����|�:��[Z�͆�*���>.��0h{qQW���],%י�z�<�C�XSp� (^P��./��;E�"t~Kr��h�#p3�/��dT��W<�YM�1'US������̓!ߠm�h�dmb����٪��dt��-�7|�e�E��l��.�P���C�q�2��<k��a�bӠ����E���&t���n�6�S����m�K�s�	�2<�f@X1V1
���`$���X*y�e륯|�K�J��{f
2t�L0�J�w����5G4�-����$����\��u,�����`�����/�mM*X�&�ðG��S��t_/�^���rZ���([�_8��������>�ژ���v��� �Zv(�!D~�i�����zp�a�h��x�i�~�"�)y	����[�*�)�A��c2�3 �t�yHo����Պ��3e�P�E�(�
�x�$8���)�񭁿+�@����X7�����'J�e���_u�}�Ђ�����H�2I�~���
55�.A�M�
���Es/F���o2��ûFt*GeUmK<4:�_~��i6�d�%f�Zׁ�kX�V�O9m�q�آWU-��~��]�U��u���^��l��p��0�&���o� 23З(�]�=w��@$_&�S�;�����V�w�ⵯ�Jt>$++e|�2�]����M^Ɇ� ~�l>����m]t��Ńf�x���)�կ�,
��Y�g5���P�c�ĺ���Z�����ck�v$A�P��Kw6D�a��4=��Lh��r�P�r�o�d�ދ��Ѣn3B>.���+/J��gT��ڪ��z�x���5��ԙ�w�\�ߤ��.�X�0�H_"5hFD�N��\6��m}7"Ks�-�g�1��6X�����U�&W���,i$4��t����#�@n!6 ��u�l����<LiwCV��t��N)�&�@��K��V��}�E~ҩHq4����4�&����W'[k�ɲ�:g�Rxk07���I��"�Կ��SK��d�<4>@�Id�D��i�z���/C_��L<)��i����z	j`�=#	+���D��*�݉X�Ô�Fc�#]hk��EJQp��H�I�<=Ζ��r/X(}i����X�f�:W= xfB�*���U�Hm6��[�����0� ��b�k��v��`Ь$��k[�S)Si�3��E&�l�kEz_��{�9�R���]����D��0;�(Ê�pf����?Ad�t�e�a�ޮl�_� ��Z�ں���ж�֊D0�R�B~����׿Oj�_�z���(!<�늃��͸���*b��GE=�0`�+�*W��Y��+�2f��Ѕdc�Y�R����M��#P�����r�F���.{_�� �4g`\���V����]1��l�*�B&`v ���P=qej�D�]c�tn��J���_��,�Sɬ7�_�2�XՄ���s|�����K�M�ÝzoTYz+f��q=���[�w��p�ų�� ��J�P�VGC��H�0b�볙��������V���5z"8��ڟ��%�z��f�ta"N�����$��u���gʓ$z��!Hk<h��wۿ�ߦNTa��SD�,���(�bBW����r�x��~�ĸ��+�_�d�4���|g�F�A� jr����j�ŋ�L��NPD(�S|�T��su����^n�p��룄V���O�y�[��;�8�=r"��['!���1��ر_6����_�"�AB��?(�;��U�x��{���@S'�[�+������u18`I�_�8X�����U��Sy&_(�t�TJ���HpT��$�L��-��-���
w%s+��z�}���ľRS��{d8Γ���L������_�D��sI9���԰}lh�)7i��#,`Ⅱ��M�Z�F�>���o>��	��(�%�����w�Ӝ[El��t=+�X`�	o���)lj+و� �>��p��:�>؇�Ǚ�z���_x��>pB�@�'����&ޗ{^��7K+p����G� �1P�*�Z�K���OV�D�L�,g�h��[����`}y�]Y�r:O�.�+����R�2�����:K�PmA�O�2*�FD�B�^��<�c�Py�P�`=�z eLFe�?��5[��z��K�&�Wx� $î��
���X���@�5�,��Ll��8��b%g�wς@e3��1�H xf;����+H��P�-Q} c���,��5+�"B� ,"R��>5Bx���0//>�"��`�xHVZ2]w N=7��5y��~�F������k�H6�T����G��ލz�{E���.�7��O��×��q��hk*}+��Sm1��q�w�z-U�G��m;i���1x��P&�g!X���y���Gw�3q�E��Ӝ�k��K>����IWL���E�9��$��t�Nk�wM%�e����R�p#���+Hm�,3>�I}�]��H9W���.�{s�)�
������	*Õ�����t�zx�z�ց� r�6������� %\����j������FpT;�^�i�l�Ŗ�4S����'˽�Y��Vd>��u! g���)���8���eg�A8��Z��O\v���W԰���H�c`�;�7iu��?�߷����g��]��Eo�N[���K"\�:dQg��*%��p��h�J/���Ή��/j��+r4�k�=�>2Cc�/�SCg����W��I�ʏd��r7��	ɉ� �e)��5����N1�exE��*,�F|�R��;[>�1B�r��O ���1��1b�����գ#�/u����k ���[e"T�>W��EƼ�K�ݕ�Wop�� S�����x�$��v�*y4#��PYR�E]�eW�l%*���A�~��>Z}=�K1�{X8�r��e@�g*��	�XGgK-V�F���_[`v�2|�[D��NCtY #��wSʉ)�?}g B�z���5LB�xn\�lrZ��ȸ2��Ccגy�d�c��8D�F���b�'%�poCj��Яˏ�\�O���#R0d��ֈ������~�ѽ��[t!��*�8^أ�Q6x�?��S��������Y$pK�:��zjQ��<KǏƸн��OUOK�b��Ւwx���E�5w>�7N!eu<m�tM$.d<a���˶Ը��#��b?���j2]ڋ��@Z�Q��FyNbr��U�Yl�G��e���c����!8S���+�F�+:��rk[��R��
�0�Qy��M�:���) �U6��&��/e>PInK+m�Ta���)�mt#�#�����j;��g��5�-�*��-�iJ��WV��zǙ�%����L�����	���L�%�]aa#��}���^��o��mn�/T8�9J�`,>^cmw4���)::��]�` n��	:�DX���Jqn㜛��6Z&t�2�p�����������I6=������<�n��;�t��ᚡ;W76֊��eԮ�o5��q��w'��THC 8�s�1�J͏�A��O�*���Ǝ2ݮ'��ɨ{Z�T��'��,l��뺻��<F��Q��C�!�b�@Dr��l�4�䡣���09�͓j��x�IH2x���f9���]`��D��Up��5�*������T����W_��5ee���"��c�̘���³,�nc�I�Ų����p��Òn��~} x��賒�|eO�8��(Ic.�;��]i#']􆱺9aT9^�yB_J�Ȩ�q��i�z�S+M�4WyJ'T��ˋ��o_�A�f�j���6Et��hM;�ǜ6Zg�3Ҝ��kx�{�4�=��'q�(,�eRY�bnn�Mn*�#�@��Y+o���p������*��&*bf@�+ן%� n����uBn`���T�S��*�o<��B�N[�@��8���>0����
�3K�@T��p``q�b�	E����/8BK\�-B�1�So�D;&=���[��d��Ҟ���t�5��\[#���><�-%�J]��W-���#����%Td��	>Z�zL�]��׌��f߷�����	����K;RP԰���!�z�þ�3�7T�i'�L�ŷwJ)э���>�J���ě41����%^���* n&���jvә?�S���Lo��aޢ֮2	�Ӌ�H2N��iuG\�^B;�i	6j��F�3E&׬�9��0Zx��}�7�\�5y
8=���e�����+�Ƞ#����o@�J�Z�r��,9��VF���Q*L$����b�F6����B{�mu�'��F.3��h�WUźy5&����~��==Wn*Y��4�m��kz�$��=o�bt���ݵ�2�P�Jɂ��8� e�_+�5z�P�:l�_)x�޳%�,V/���6
�Qn�kaSi�1X5���]5��]�pE�������5B�����L�}��h�m�}��P5���u:�S�/{�%/��W20a����~�tTw�a,��p]�3޶\*IZ��c@OǬ�"j���d���g'�OYU4�&����h@��������}�H�t���X��k�(a0sz5?���iX� ==����S����;��v\�^ߞ�>�9�!����P9^�L�DoK��RVʌ�[GzW��%���5����U/m�:U
�08�SѤ��f7�j~J/r�O�/��yk��]�=7�_M� �+˄�>��-{��������TpwR�R�u��.�8���#8n�U�P���]�]�� `��r�O?���ثJ.�_,,�l�D|��9oY�U.��̸��ΑS��݇�9���~��h�ۖ�^~>俉ij�$�CCU�X���'�%��v:M���� 8=}&;�(8��5{$���<�)t��ZJ�S��j��Q݊�*���aR}�܈�}8��L}����#��:��(��D�o's�42L��XW�~�H{n]=���0�����\�@B�H�Ca.��h�ۀ����iAqȒ� (�3�z-ö�ȶfP]��ʓZ!��4�e��;P�b�����1A�B��XA�CpE"wq�����<��qzG^�Ȥ��q��7�4��8�9�����2�D��0禾��|��|��O^z�d��D{[����E�orM�.�K�d{��y5�d��ĝ���nīF��2"��BSe�}޵�+�S��]��Q6b��L����^����\P	����`��f�x	��U怢��Ş3�@�
�$Gw�o���}��0��<ح��j���KDa!��e�Q�z��������V�7���{�qb��+�L�zt�>������evx��k�d�0	�}TE.����eޢ��,D�-�ż�����*(iݷ���&��k
����V7&qb���d,�A�w�e������l�\'B�k�=
}`j�y�nm�Z?0��Y�ӐS9��Oߋ�*E0 {�������A���b}>�ܣ����;ŕI �W}BV�5�>���J/Q 0׷����p�E'��1� ZXGY�v�,S��5A��>&�����(�z�F>g|buzq-ru�^ED#���l��o>�����<���0��nMmSO��,��M�r�$�}�{CVj9�`(,M��e��5+,^g#\��ߩ�d�D�
�:�мA��6\m`mٸ�ٔa�`U��_W�6�Ӄ�h�RΗ�@v��J�4i0�vδ����&�g>�
�W�;���҆9��H�N�Uρ�����yI�W&tاT�$�#��Q.'�W���x˫�MR;����U2�P�VTY�N0Ci #�Ef������+�y���G�5�ML_Ϙ��8X`JyT�䥪'EH��4C� fN~s� { �;>��h
�R�Bt��s+�4�y�M�	�
����7�S������۟1��}����01�ED���_ϟf4�߭�����T���}��oؒLrJ�=Dfp�\Q�
��''�qz�ַ5G&d�9s��G���6H�
���Nk{��(z�T���)�xv���XZ���H�"��;����H$��:���JR�&G��E[�߬�,�Mˇ�IڜT�%8����>`��NT�t����0�/�8/�3��4� �����v�Y�.<��:}ؾ��G�K4Uzh�ʉ%#��� r�Or,�s[/@��i�٩�:+��[f口ф'�L*{K�E� �ʮ��+�����B���UĠk(Y��O�;ϳ`14�b����\�!_��� ������l3����qv��z@��)np��O*�@��	�F�Z�[��3�ߵ���ًk/��M�+\2�7f��'L[� ҫ�]���?_�	��)��S)c\Q�}M��R�8*	��mzi�z�N+�1���B�N�V|P�k�ǩE�3���'"MV 񗭈뮶�Gߧ��YZ��~"�����; �e^�Rk�t)���6.���@=�PK
�do�{q]��.*븙~� �$�#��9�Yx�(_�K�b�TΪH��է��������O`s%��0^�H��n��Yh'�EҬ�ғ�T��62�����.w�a������r%��5*�9���ַ��gҍ��Pt#�8��]ݑ����S�W��j�^0{���<J_%����΢�`Κ�̔�Cg��M'�=M2�	O��8o�:��Z�(��H-|����h �q"����1<e��j�Q���2R`z��c�0[�0�8��N�pU-Q���B�VE�3;�h&s�LM��SSC8�~Wy�+ץl ik�)�%ԍQ�A����;o�t3�
S�$�$ˡEt/l[|��p�?�����ĽL:�E��G��m"������ٖu��ݕ�s��8;1�#Ĵ�m
=���~����Z���H�Y:E�o�ק��������3$��q�*�Z%M�]#����:S��dwZд.y�]z�Y���z�
�n���3gtռ]�?�_���/�C�gܲ��>qY=N�AW�Ir��>�8"!��Ǿf\YO5�x���@��2!e%��ֻa������)���w�R��b s��>1��c��p7{�5륟H�O(|QM>ZU�M��<�L5ޝgQ�$��G�g8��a��ƍ��"�b� T0�3���vgZ��3�9�e���(Q�.M-r�\��
��bG<QͻB�Ar��4�z�����-*��L��v�Jk�/X�IP�\1�+�ԭ7X8��6���pI&�/F9���&���!@�u�#���� X�|#��H�s���6��w�`.-��hF�M-B��%_����&ȩ3c2Q�8mb#����[�\M;��$
P���\�({Q5��I��.7��0)�|��S@�1�eȾ�KJ�+�����7!�X.$yQ�X�t��WE}���B�V�h�Ȍ��7��(]դNV�nbW݃�!���zAE�.4�'g��/hy�9�C�`k�]�,�t��?����!z�4���=�н�N�Q��l����7��w�(~ۍp-��T��c#'�8��kc�~����s �Nf����� �x��2���k�r@( ��pZ5��F�����S��R]��4v�%A�h��������
���	�@�_�{�$U(yԷ�ϙ;��̛DI�:��D}�\lk�b]�Ftw���m}#R�d*S+�!�th�^������u��~�ʇ�n�75>U�	�?]L�F�'PA��u�c��F[󥱺�/4|i��M�p���y¿��z֪�!�!���>���6��?��q����w���=u�Y�W������b@�<���<aX�|��!#��2����N�A����2���UVX7�I*B��ʑ�<��j�u�kҧ���������U���@, �������c�E~Br�! Ѷ�����ӏ����(�A`Isw�eI�~���h=d���xB��X͈(��G��H;��o�T��P�p �>y����uL�7����Y�vw�)N��+z��C�c��a��u���ǡ�/|WFA"�P� ��rІ<t��kQ� �P=���{ �_�z�s�b{��V������L�_T�l��rc�E{5��)��Pr�٫H��Q-q�z�����tү!���X��N<ΙL�%��D��9��Q-� �gM�Q���w����n,�1�ٲ��,��V��N)prU2f���o�����j�D�w"�5��2�d��S���9��|K��ƺ>���?YO���]G���c��� ���P5�ﻱl����ќ��J�(t��rܹaOQ]�n1�vy��рS�Zp�K�0/P���y�㆚e@b��G���9v����� u�ߍ�;J����C��	���g�}�=�_1t�]��>�h����Rh���WO��!uY� ��{�D��C�-�ox����� >'�AO1ú�	퐼�.��rBW�5�<��a�1��\k<��C.�y�b���̥3����A�&��K���;���cԩ��cllE��-�g�~�L.q�ѵ�U�-��q]� -�q�;+ab��A벓� �{G]"�1siV�eg�QEW�̭@g_W��d^�
��g�Ű�X��~�f0OG���d�
9؎���+��ᱬL�%�Ub�o���v�0�	��Ђ�۶C����f漄/z���ur����O��SAĺË�/�, �^��7EoML	KmD҉�Ȣ!�}l��h�����Wu?��ݨd�A-r��x SR'�W^_��\C�HL*h�Rޗ����Њ[��0�7\�9���j�0_��jp����G�w��)}�m��g��[���@�dɯ��lC�|k�7�ȸ�jN�~�R�0��l�>%�/�ÔҲ���=#�=���f?�PbI0��Xa�?����M�)�f^S�����2�O$g�d+�>5m0��ZP�ʬXL�xq^� �_�#TF�ޘ΍8�o��\���"F�t�}�F�u��-
CqQN<���nܯ��~�I��+M��Q�B9Wz��
���ْ�k4kc�)`���D��q�[H��M��?�0f@r�}&`��QG�˯���5�@-���7;"�u�ٖ���4��V���;h�� �h��ī��ⴈ���c婩ƫJ��A��P��l����uMh��D��74��5�)l[Q�E�Ӝx�c1BY��>Ґ�D���4�X��x��ZO���I>����5�}���l���_����.���㪺0	�,����B���
q��&��#qqX�e��Ts�P�6����J�i��O�a,Q_�b�K��;'OѢ�5�{���{�B�-�8al:�v6J0%���l��EXz��p���:�����M��|�f���<
:94ۂ_Ǳq�&�KY^ՠt��ʽ�����1���ȃ���5H
�����#��ݻƫK��|�*�r�p͇E�ePh�F���_c�6,-t�^t^\~¬S�Js��� g�ŧ�?Ǣu�^�F�}��6�����Y�X��ǎLЂ�!p�����r��=!�5Wy��_���� ��?�+�٫����P�r�r��ڋg,�g5�|�zm���18w�<���oDE��oqb�>4��3f�삽�h�8%�i��S���A�Vx�:��^�b����qW%ΐ���叜ψ�'�Xd���<Rp4`���`�� �꤉�a�aR������ix?w�`{n���7�)���0AqENL[z�1]L+'�2V)g��b�ߜV�9�x	��f�}���Tq]WIL�.�r�"A̋����.+Y|�.��(z�lqU�J���o�<�0T��b�W�48�mW��rhC+������W4�?Bb���v�d\��5
J=�A$ĸ��eQ���X��_z	��P�������֌�����EQ���BL=��*�az�#lik5��W�sµW��}p��Re���|m��ļ�z�?�#M1\���6[b����8�υTt�)������2:uC�P@�5��1�t��g ��(�E��y��B+4gɀ ��ϳGx�0ĭ�jE���9%��c�Scώ6?f(ju玂j�&�|�x��I��6�Y�:�IxN�VM��I��sD��2��H��A���08ŪS/K�
�B��3f6�s!��n�5�G]V�����Ќ-�5�E�a";��p���b2���s�jz�̻_EfX�x�t.k��N&���a��� Ш�=;w�ٿU�g���f��l�Ö�g��uMu�p  i�J�1v�Г���x�KŘb4��mB�irq�|�#~�/�����!�叔���oLm'�!�i�p�NX�A��G��
���\��g(��q�w��v��kF ����p��	�ïF�x��U�<�h&�xYX��Gq�	���EF1�� 6��\"��UK*���������%3���ZGI��OQ�J��-���h�b����P��jN����w@��h�*���Ӧ�{��u��J�KML�^更:��^�+��dv�ւNt$Հ^�e~�5a�r<��+x�IQ�M�~�B�w�2�ƛ��G�ǌ���G�gͅ�����N]}�E��K�f��}��~m��� ����
U�|	��e5�5:��l:a��sEi�[}(�Ѣ�������<�hr.�U+R���?�J�C�Zl��!��U[�\�y��v�j��M1y�w)��!����	�'&+��9;c����M8�����5����Բ�j�ŝ/�0L�S���d�l�ecD�s�<8}�oŐ�΁Fl��4M���B�,��	�L�Ԁ�9,D�A҉����9f��W��5�@����s�£��3k[�)���:��\�a)���W�wsP�78q��i7Se���6�!���W&�
:���#^���&�����Sfv��#?���ʺ��>Ku��5�*/{��6D2���F����ߏb����$�c>��[���9�]��w��<^��o�I�Ǫ,V)^n����j�th�f�۰��uf������"�~�,9���u�BF �6��a.iĢW�*B�T|���,�����N ʊ(����_+&���'%B��;F�@��2C�΂��V+��+��Y�+#SaD��Gĺ0��$qր�혳ghK$f�{����b����w�c��G������1h�L�E��GP�l=e�<�@g�0���WXɯ�EL
e��5pcY!��b�=êz�U��xr���݀LD�Fk��\6Jd|���ż޽�����:d^�F�����P�o���A)���Ԗ�A���)?[ ;]VBR��L%��}s�-�4�k6�B� ��U��$�i��|RȊ��e��y�~ڪ�����`������O�	]��؆~����u��@���T�o�Ƙ|Tf�~��Z�-@�e�"�;�
��.�~x%e��eU�']���D�*,+�f�̖_�Z*�؏E�&��G��� `��8Mj�Ǘ�z>/��p���|k�uaGv4���}1�\
�ej7�"ŲBX��^	l����#��-��;�L�a¯g󕾴���� ��ak�e��噸��N�|&���u��W�x�۴L�MK/�%��]_�O�#����%��c�x5STO�BrHԅ\۶�1�$��8����ׁ���e�-�D�U��(?�����@�@���,��v�'?Fo�����K�>�do)���&���)��^)��A�M�FN��H����	OI�,��&��ѡe���l("��A����уJ�m�4��&=�[����c��&(��9�C8�!rZ���O��y�ٱ����:��ofCF���^#����
��W:��D1��䵭aqÒ S�5_�s�[��YH��e�CT(A˶�`L�s=��3�7W3�G1�H��Jƽ�H��c��^e���c��5&J�ZՑo[F}S: ��WH�h�KU�f�!�[ﾨ}K^eoB�a�p<�*�Z]�`���?�5Ag�S&��v'��L���H�i�(T�uJj��D5e���,w�Y�Q�)a{�����̼����o%��TP�t���q^Ś�~��}��F9��\I����R��6�A�kp.Fu�T��*�0�ƸR�m0�I�-$h�h�y���f��@o��Y���Q:;:~��k�*x3S�V�������Y��IKpc�<��*��>%
�$���|!DZ���	z�?�m]ugL?�M�Ъb�遊�oh�t�0������U/��om\�
V���I��r��6ܰ�_�Jl����k9���lft�{1k�a��Ǆ�;�?�w��g�ꓙ��AcT�8�.�99��uz�2@�|[(����p:+���*�߽���	��R-�8��;��>��
�[�kI�I������8���`1C���t^i�D�S8
ɿ��U�cX�V��c�S�q��5��U��D4횲M4p2Ħ"5����D���
��=����J��J��𧚄a�TQ�G��c6���n����q�;:qKY�吺��W?4�w�q�����M*����mY��[ ��� ��-���of���i��C2; 6C؄�3`ࠥꒁrrD��5ʐ��ӡ)\�Fk�Y����	��r����/�6s3�X`����T��.G7CƏ8���&���Yl��鲾�)�լ	.�ɉ��7�_�%,�F�÷����!�@�V��R���b7�<,�ke������	-��a0r� �]s��`�M�H��H��
K��f�*��B�q���7�k��7��ڲ{�H��J�Q��b'I��eR,�Iz_H_i~��x�]�vwO:lg�:q8���/��!�����vdj2�[��cZ�*��{J�t�|������o�a�M�9tv�p<�՗:ǥX=2������l\ҸVb��T
��ͻ$���}��̿k�w̰��-��sY=���1���F��AjK���fB�_\!�0�%a���ҟ	m6`�(E�QH~<xnб������a�[�c��$��@��.�j����n���R:���}L�ۀ���v����\�z��Jv�J�Ocb�M�����CE�O̳�c����Zd�X ��"�����(�Fe kJ���w��L�5[`�5��C�A�絙a9� �G���N�m�$Q�f�8�)����o���->�:
'� �nq_ZH�{�UpS㺱��b�
���ҟh�?:���e�񑟧��h���=��}B���,�XdF�����h�a7�jN�M�g�t�}b�7Ѕ�_�����`� i=�-�i��nix�����D�ӣ�H}Mzv�m��:2�)��؃�<m� ����d�"�a��ڇ1Nh9���Mn�^xB���pf"���R͘$����7��T�!�Q�X?Cī�}g{�yA��������ܑ\i�a�������S�L2�Ɩ���������ܨ�~��%��8�(����ݍ��$�^5�L�q�q�q������vm�nr���t`��rUI�Pr�8� gpUr#E�1E+�8;�=��g�!P�>;D������t>�%���Nd�������mz���lS8�߳������Ff�	�ܽ�3=�bX_��k�'n��Lj�G��Q��z3�H1 �옷�<��}�;��dȕs�J(N8�J=Hm�/>ZKh�2Y��NCk�8]��)�-a�<�T�T��|:�L28:��!�#��֝��)78�cYv��1�1�D��8�9��� �)�Ce� 8�M���G��� ?Ҽԕ��U�������]��I����a`E���[��e���6�k��ǹ3���]X�#�q�E(�6���g�,�\f�D�y�r�x�\+t}��s�����Xh䟇ǡ��<�D���V��+˩{������	��u��{6�I��Â<t����"�T`а@ep5�j��E�E4��O;�$琽d�ǕM
6���u�+k��	|�ٜ�0
��G�ZR���W{6�O9�˵������u\�5tg�!���K�i9̳s�8�}�����kx�Ld�YT[I�:Z莂4��W�
)Ą����a�%j�]һ��Hl�R��l.�X�#$
�1ʎ��O�P9�RmY�JHVj��)�#�J}5�a��S����M��������M�{��N��M��Ct!����S|�x�i� �r����L2�T�7P�L5���'���f�K=�cD4bvA�Y��(�^��ߊ���c�~��-��P���	���SxACO��i��7NF�� o����+���/:�A��	���x�'t�Z�Bz��W!`Sf�_4�D k��$����h�׳~3��I"]���xeG�Q�=��O~i0�y���UQHA�<sq�9pL��D�2���Jݗz3�!��U���)N/_����[�^#0��[�V�5�;�cgI(�m!%��	�%~V��5��^o7��ɟ�	J��|&�!&�Nc(=����81%P�u5;T��ؤ�B�3^�U�F!���6>2Į�
��w0@4Y2� Rk ��R�')%�-P�cQ����S�3Y��$]��b�<��t5��B�����5���2P[���6�!w����H�d%p���`�*�+��	���Vy�]|c1��f����L�.�ٔ��5�|�[\h�_�$C3���{q����{toC�N�43����d�g�"�^=���Ji�<�f�k)���E�K�?�<&�O�zR�����{�P�@N�)�*ם�%�62a�C:��ŭl.&�'vzHf�_�vO�yV��"��?�n�Fg���R+�
	w#�9�P�h22;������>S�P�op�{Y0� J4��u�5م#�N�~aY�8z4���Hi<�}&�G[w�4I 'ra?,L�}�l�^>u1�p�S)h��^�������:!j��7o&�o��3�B��қi6�#��Xqюe1\����L�Hl��2�JM7�.�4Z%[�Giٌ�E�b���ٻ��&z!4Y�1dԻ�c0���D�[c��J�[p�XN#tv]�"
��67���A�~M����X��u[c;���0@�G�E'k,�\�o�a#.�b��d�Ą�goOW$pe��A�g� Q���d��ԹC@#y@�o��[���L�_e��{��#&Ef�].��7`�hL�&n��!�PF���� �V��������"�q�<�tר"���t��:$GNL7 מB\ �j�P�2���7��m6
�SR��u�!+��S�,�(z�1�Ӑ��OR�2��?3�2�����a���c�Џ����.���e��&�3�AA�*γ�����}X�H rl�l��:rqNL}_�{�e���~Gb�Y��:�!2��H/��h7�'��|Q�U%�)���0��©�6,����Tv�ϸٽ�C�hO�G����`&�:��.�[Av���5��Y�Lޢ��)�r�q�_�*K.�Z�e���K,M�=�qԪ{�W��i������lz>���\qc~M�1��[�,F��LF��/)9E-i3��N���*�>)۽ ���~-	W�S,\��	�`;��\��iF�D�d�1o�X��RP�j��}r1M/�l!hQ�ho�g �[=Sl����_����Px��r^55Rn&!&8v�PZЕB�����t�<��)o�IDbnlq�g���Ou��$���V�Q\x���d���/!+yF�j���5W:�0� (�~/���ӄvC]E�tg�ƹ��#0h��w`X%��a�˳Җ9+���F�>A<I��9��\RU�^V�qX��_2q쁟�Rs�:����7�����rQ�n�� ��K�Ӄ: 숦 ��F�b����
��6�Z��(�$��ө۷zZ���� �dǻZ��4_c�\n��C��j i�椠����=�2X�`��wܤ)o&�B���'!��OǢ�9"������||�� �咤)j���H�`w�!��}Ҕu�N�HpjD}��,�6 �2����p�݌%O��v��}�k��~)���
�$̮���%����MF���8�{����wL�p�sOR�>���3�����z��V-J($_���T*r��T�ÌRρ��i�#Z#���΁���ę�n��1���IO���� 6[��h��M�D��+Or�ځəY���+7FKq��6��L�M�;�5�(`,mrY�pm�~˙���T8��.�do��|��w�n��^�85HA�7��Z"��N��+����7�d�B#���EE
E��0�Q���3]Xͷ��&�-�s��+y�l����9Ş����\�X�b<2��(�� u���J	��-���҇K���|��Hx�9oW�Q�])o�M�7(��-���s٧6�`�ݳ ���E��G˯t%�i�3M��r.7Bb�#�Ȁ��g�nb�O�ܝ��>�n��ߚʧ�w9��[�.�f&��	y4���ܢ�D�)�<"O����Է,F����w֡(�"���X���������I��]���(�q:#���k��NO�_fV��3$�3�6�<3‟�-&�)aF�a�2�]�%B��4ߝ����&���:5|�h�I�>��=�F
y��$EP_�~���\͊m�N#B,�;�g8���iS���c΃ D��.����nX�?��]��ݠ�P�D�v��Cx�|YH7��$���GCVo��{�͋���;��T0�{/��La�%l�='�bƋ`f��t��v:�����d�3m�Agww6٪�
�t2cP`���P�h�Q��I947w#Ђɯ7)�݁��L�[�eb^�;�#9��5��٪�u�k�_
��V��x��$�����R�������	AT��=�%_弯e��}0�M�=�;��7�Q�/�D�M$�HR�G,��������i��X�8�r\���M���@䗔�;�*��� á����\��n�a����B��qlO�� wgI$a�!��f�Ѻ[V7��ɼSp:	��M����J)�iP$Uo��/J	Ü\/��ޑ����rYD,�䦲]�F N��᎒��0�	���^��o��_*���v�<p�B	%��1@j���elTt ���c$_��No�T8��}Iz�̈́��M�����E�:N^��6j���M
��/���_� ;t�?pO"�|�ډ�_�,�y�m�����}w�4��J~#�/.1�c?�n�Pޘň�Xf�?�6HWH&��Ft��!X�u�SHL���SO��+�Z���fyw���( R��&�q���ś?���v�o�7�0�ͻ�%W��n������p�e�`�(�"��M��O3�}�2�E�v����vF�� pYNsT���"���B���Sκ����|$l5ݺ�\j�ti�~�_�6��|Ƀ`���Y��ՅƯ����M�7F0�m�	�b�ھ\�e6K"TDW1�h�����[�����-��o�s� T#�b���]g���CQ�7�+����?���];�̤}o.ߓI��?51~p!"�ދ�<��us���;@xt�赵����%k����8Fz٠�lT�
+!���;���\.i��\�ʉ.. ��q>��|� e޴͹A*�N�5�Ba�Z[N;���!R��	��hG���� >�X����k��E��uQX�99��:�7Q�bUT��W�gN�����R�.��ڨ#Nc�6��Х8s�:�N[�鿽R=d��qP���C�V)M<n�ȆƜ9�-Ʃr�k�G��C�S�H]]��K�  �Y�<�՞���Njq��o��뭜UH
�e�0�?t���?�\�����U�T�օ��?v+�J�u��90Ӿ}9r���aGQ���gN���.-�R�\��<�Y���q�U��g��/�˕R)c�gm�flː�g)�]"5�I�Ci��#� �:1�ᛕ�m�6�w�w�`�22�oxw�q����@�{x��r� WA:�gzT>�j�>7�Z���+��U1�{�|���ȋ���N�
�?,���a0�����@F���$Q9��(��`j~"El�	ҩ�߼;�r�ޑU-�9N�R��i|Q�"��?�N�:���q��6^�$�׭2DV�^��z}�⽙
OS1��ZK��:�a�
,���w�fͮ�m��rܾ(��%��5#���y�� �揁gg9��?24�%ud4�	�J�h����D��;��R���׾v�8��8��gTh�;@��0wt�U�7�3D��i���9�p\����N�!��c�p�1O��t�T�?cu�0Y �t'/�I@ۂ��	1�m9��]���dۢ���R��@(̿c�K��(?��W�$�������3�M�x��9>]�!]r�*� �SQ�Ҏ�PǤ�_^oDT߃�^}���o0��"ҁ`;/�@���zNl�}�B��W2v��-���U�6�r�2re)|q\��87R��-2=D��Y|�œ�:(u�]�V�s��Tt�ްU���Њ.C�ܑ'p�2���H�	�q7�!��l�6��g�=7Wu���|����v���͕��.?Y���d��4��w���I�Q�kM�"og���[;�F��۠X499�Ty�AA$�j+��}�Z��v�8�<��=�:�5k+9�S�xj�tmP��uNfx�\-*� �v�x�	fq[P_��d<�=�iH&����d]��l�_S'�����\�!�M�E�ae�/hR<�&G���b<Z�uw�O�5Ro�<'������ �v/ξ�5��<�Ѓ���}�my���,F=��X����c�i磙|`=�
�7����ÊEyԣ�,z�5�6[���wT�hnJ���@L%ZC�R2�"}���>]��j�)M�#j$�h+�կ�|���(���U^+���<�s��kA4�^:]8����y7���(�c� ���w	�D&1�E�T����c�1�ƕ��|�u��)�����ig$x7(K�>�`���u�Q1Z��zH�%m�y�ɪ�Ւdy�U����f+�'�|��l�zL�Y�+<�8�l�`Q�.FV4.�b��;�9�r�x��ֱ�E�����ْ�k���rt,l�A�$�V#"�gzv�Kω)P"l�4���:M�J��!6�)GD�P�݃��u]'����"%ņY㲙��M��Q���D�����$r����ϑ�/3��Z����샂�,Д*�&h���p��*m.$��)�(t�<��%��M�Ns���A\��OM2����&�[=�0.g��Ö~\E����º�|8P�\�_��4[
\�jM�O���k�F7�H´O0�j�N������r�Ũ��e8i���^��}F}5Axx��Y��6�/�b�'�{�i��==H��H���}��Y><��W;���j���1%q�K�;�E�<�O�TG:dG&Ր�l��Q�������A�1|*^;���icm��(�<+�7E�`>	ҳ�W�����*�Y�����?�@xl�f"�W���޺��`w�wA ���'F��2.`���ٞW+���#�!e[�)�۷��W����w��KL��ʱ|noC6�"٣g7*a�]�U����C���4 ��t҆�1*�����zjx7t��H��Aɩ2��L�v�"J�?���tS��]�`��љ��M�$P�[��e~�;?Z�T�.
;S��7�\�:˶|���(uO���D)3j�]���١�A�^�>������ܢ������!+ZkP�)��7A^�<F;��̚=S��v��}�����lY�:��[�j�nݰe9�i�5�kE�������Q�	�QS ��LO�
˖������_X�g�z���>�UG~��pGi��7Nak�y81��%�,��<�c��C�o1+⪄V�4~zB��БP�H97!�/
@v���,��QC%j���%v��㕣�Q{A�8����Qq��!�ƥ�"A���\W 6�єӌ�+?���^���K����s��P��4���Ï���4�ɚ�|ҧ΀����,^5�؜��Ms���_��B�1��D���Mݭ�G�:�*eX6�6^���̵��@0��cG#cNp;]2��t���a���u�ݭ�4�+�f��*��)Z��Tee�/����-�x��R��V�ΐ7t���V�KzTo��¾L�c}�\��8:	Ag�}��@�qY��{�/T���n��9@K�`Mg���M�*��]ߍ�S>�?3>�����.�~tb�����\E��܇8�~"���+Z�Y�q�< )G�O1*tS`�쏳*륩c��2��͢�>��L���pQ�l@P"6X�T:����Fh�ҫ��:���b)~/.��FzwU3����[b�ճ�W�0"���jC<�M)φ�(L�ʠ�o
�OP����
�It�2�V1����[>�ZG2��yfCg�엓��z������ �������o�Aw�6�0����u�{��BV�����٠!������8{�#��O�v)��]�6qm�yݛ)�"�j��y�
��ʸ�N������`��6׾2��3	'o/��[5(\3����n��dIm�)ox&h	�hC(w�|�8S�X5��oJ�%L{��M�\f���3��+,>�r�	Z��}k���Wo�B+z��S���e��zx4���[[2!�@�G�p�YȬ�1�7��(������k���X|����	�#.q�ޠ}
R*v�S��;�R��H�>se"=>;܃�X'��g\��v=�Nm(̯�����8@��ڷ Cj�������X� ��\o �c��DN���$r��:��l��ϔ1/��1���<>�� ��3V����$��TMP�e3f�?�Q/��怃�E���pޫ��˲-$��:��>b�+���W���ߝ��+�S���I�KO��K�-"/�^�U7��E�1�r��������G�n"�L�.�m�|����jc�����{�R�M����k0%k<n}ֲ杦�QQ��u���������By�>�CE����^�d�[4l �
C���n&Q)~ͫ�䦠B7��#���մ) y�N[��G5�W�lL 4��X����~}a������V��l�>D�f�C�L�93lF��./"rp,ȇ�.g�y��e���ݹ���V��v Z��I�@W1���]vpYk��+�V���Y˩�>}y�������ΐ��s��5?�v �L�;ˌ!�n��x������M������IR���I�����0n46�6��,�[�1��H'��4e]t1
6���L��~Ch
qnR��U[\ań�j�N���=wi�BΆ ��2j+c.kԈ&7 �f5��
F�J ��m���x���#��j�)8(59���wh[��M�����@��W��G�l�.�K[�=��Þ���0)�=�(�<�K�a���c�
S�ٯ�]��g��ֽ�ݜ�A�'#}��7v2&��{@(����̅�t(�Z�|�{��('�ν�����詭.�}����=�$bOH�܌�?�fj���` T;�V���ʬ������Vcr&��Z���[o���'ft��.�v�g]�Z����kT��Q�=�̦��ءGt|�n��1Y�QS�`4*Q�	�;Et!пe��$���R��.5�*��罤��'?��Q����\n�th�f/�F�*�H�	kG�<�UW��J����%��n��ED}
��i`���$i����L�KyG�rU����OU�Hx�R��Xp���L�8tjQ:��}�斘"��Y��㥲iF�X�-}}/���H�]_$��[�yrƗ^r�g��:j1�
K���9S�����Wܥ�� 4����G�4���f�U�����:����~&���bUp�@Am�"BZuܚ�~
����s��(���X��(�
��Y�S7��=�n�j~�o*�gr5}s�tq�C���bLC��@��l򚰱Dޗ�6�x<Ԛ�/��������Si˺E��&p�3<�ۆ_�HT��pM��s=h��Cz��tP���$_��R��	G�7��ݷ���^��u �t��k �����`"sd]�43)2T���6����)�Ոy�mY��~ӊ��Њ�J�5����e���1��+f�.ę���EP��
y��}Q���)u&5�hk��;��?f����5�M�PHK��Ob� ���L1�}j��I��oT��(��a�r,6N9���GiI���Q7�^8���QjO�F�1|6v�ו�/ռ�@�;���z�� �%���T(N\rY�-E��Ք3o���}�}k�������s�L��պ�i���S�`i��>�W_}�C �x�xA ����ֿ7�]�K�{m+LcR�(ܤy� X����[�������v�\���Mq�U׻����S��>H�� kaN��;3��:3���cI��D�p~��w��C�)Yt_�}�G��W���.j�6Z��4��{�,�=�<�L��O�l��\����Zp�K �� D��#dӘ��'*��t[�4�Q*9���D�U��~�}��w�P���s \�7�nuan��T�J5���?
�'���a����+a��\1Y`�.U�6q�m}^�Ήg)�6�@�X�vA���WI|�Ys�6�Q�2iI������4�&������F�<�>�>��/���Q����� �<��*�}uh���Ţ�b<Po�~��I����b#w"��,� pJ�r�b�����̞{�5SC
�׽s�/<"��Ff?lK���]Â�G���g�G,ڇl�Q˄u�%0�m־���'���F6�?]r�tBP�L��=�������<�,cdhER3��+�!�<9��t�gӉ/vJn�;E��=�a6 <�|5>���^��&���D�~��w����K�X�s��MX�e9J��P��Y�Gli�Gj��X��z-ܜ��B��G�N(]�;��"j�7H�<c����[�j=��Fc��v��@_0���;`ri���*��v��Z @��K[��weq��N<�W{R3���p�h`r�r���z塒�t;��'�o�'���9I"79һ�WY0k����ʕ�p=���k�n����ޕ��?^�?�I�������g]$Ě���׸�_K� 	��)J�Ae�,�H!C�cY`��#��6����`H�_�X�-ΣbD�t����T�)���r£-<���dac�am�y	"�4�7���xK�m����ZQr֕����y#�VdD�"7j��n�kdBPq���K��k	7�h�qbX�D���.Կ@"I^�!%��V����_��h-���0�ā& ���^&�&9���4��Q����V�d�VL���T2SB���r6<�^�R�D���
u~���@KQ�F8?9�aC��K�Q����Sl�ĝ����s�4���U������E���_w�d���F���z�^m���S��ŉx�T�ڝz��M��x������xYƉ����]xtJ��1fҘ-v��q�?����+�|���Q�Q�vC���15Ve �b�/�����P!��f�5,����
��<�l�[�p��0ځ-�Ki����N~C����\�Xg
����\��3tͮ4nDM"��ڝC��%��t��7r毅�w��T���A������}
���U����GVq���u�nD#���O��]
�	-.��~��d�?8I��66��@��E�|Gi�| �b�,�<iͲ�8$�QN�	Ϭ�ϣ�^:��-�w�k�q�:\sm�^	����ܠu�&�|�	q]K^�ƹ0���?I?4("7{�O�Td�t�{�3
���vj�r�N�^�U�N�˰��?ʤ�W@|tf�����5��/F�řxM�$��pi܌<lj��3�=i�Q�X1�L�L�%9�t�hP%<��A�ц
׵�@B�+�r�ʜ>�P��_b�&Ŏ�R�y�?�F��2�]}K&��ks���86~	��%���`n��[�]�+Gg�M�	�	jD0	(rE �:�	WbwӴQi+�`�@�`��zM��������0N;��!�jI���:�x��t���/�rw1��턭e����5W1�"�ZiU`��qC2]�X���C�f pk���t���N�����)��m=8p!^b7e�t�lʨ�5e�9�M�K?�q�2�.�]-��̱U|0hh��ztJ�:H�]e�Q�tAn���WV��Q,&���E6�E�'6C7�[˴����KdA^o�!꼝�	�!�y�!����j�x���\�o�������͉���L���=fTN[;�Q��B�Ԫ )z���ҷ��ʞa)��m�gC_��WD#����T�w	ǝU�z��J���_%_I�/y�
	������GR�8��(_,�7�
-
'����f:o�/���\x�R�a�.�f�^���v�oH���l�Ȳ'����r��������mƭ/�F+=.��P��XS�*"��O��Q�ԓ )ι+���򼭬.21��-'�pdo��'퐿��U�����L7�J�W�I��O�{���Ʊٵ��/�>��X!��?E&��R���2v-������:��Dk��I�5<l4����S7�_>m���laGP��=6�x
�&֊,����n��Z��b���K�9I��W��->g�r����y��yL��s�:э�D�K��e3�Z����$�f,T�He��=�����6.���]s��[����������L�~a;��a2���cdmp�"3!�y��a�AŕZܶ�-��M�@���87�mnj��Ipf仁�i�M�����pe�[�E��L�_�dck�N�\��	'���Ů=���V�K�&Ӂ���<:_�k!�K�eǱi�0X�����V%�hK*�>����Ո�+��M샏T������O�(������t5���/���6��$��zA3��)���H�����b���]�eh��iYaä��6]8re��]D�8��T�j*s�e/�M��G]����t��,#���"��A��Lب�l`�O{C�]>�i*�wwl�T&Z��}�>ly��Ƴ��i6΃F�! �u��`}�f�;N���?b���Ĳ�������r9(�������"�*k�bu����Qi�oR��W����n��I@V�;�-{z��+Z�e�'��IE�u��	�a������t��x���MpVt��� �l�����ƱF��7�X.IHLtԑ���뻨����-@	f� �7rn���M��a���,9I�l9�^lL�Z�5d��p�b�B���|�Q˕١��3���qO0�+�?�{#�~��h�H�#��ќ�ܕg�920�.���mb�m����2c��fഛ����b:P�: h�Jh�u��Ӄ4��[Kz����#�a�V'�h�0����u�Ϡ��W��BH \)�4�:#j�'�R9|��N��ɥo/��Ez2�QH��>�Dr2\6Zw�;�\$�3������2Օ�v��}���Q����T�rm����qI��Jfw^�,Ƞ,��o�	�q��m���-�>$)��7��P?�����~�"䭌
��q��.{:�%�~'�B�:��2M�eI�m3N���s 5~a�[��G&�\�Y{���i��XȨ�E���?�?+�7c����!��ٖsg����PQ2��)$��{)8��"�P=�g��g�a�����%R�/j,�9
��#m/tn�9ԓk�)��Ta�1k�kJ�i�7n�Zno�Z�~��Ct�9l�[�_Y�Lo(�ש�^Z�_`>�����s�F�3���#�j��@�ml��@Ę��/������s�$%FH�V�';<�����YVħI#8ek�Ɏѽ>}�����5i�}�zu�\]�rF�E6}�v~yqVw�}��m~�1�4{T�4 ��Yk� �',%�)�i�Y��⪤P]k0���p��=U��(�%���"C.�X���\W�'#����p�nk�Z�l
A햂���m��ugXu>���z���@A���YF^��ǰ��IyYPc3����j���MǇ?^Q��x@�>.`��Z���:'���0��~�Mv="1��+A�@G���ԫt�v\��#G��d�e�17.;��~"p�S�c���; �㌯y��|jR*�}�
�eT�����~��w��'�1H��`�WKca>Qg����{�5)�
�+>k�7�R���F��+�)i|���I�JpX&ػ���H�͟��[KC@|ܢ���9|D=�M9fH;5�G�~\��l��^A��}�SɑW��<+�����Z����ѷ�9���%m��Ap�g���V�a���a!���T��{��J���K�j�%���6��ynO��;��D&U�$`���;$0Z�{����Ê�)���yJ��}��W�F��M���w�V�C>1�0O�V�f����Aw�MJ���/�{uN^K���N�����=���E�L6ڽON(^�����ԵVYg<Hr�q`�J|�M-e�~vЩV�w��Q�N���
�3x���+q�*��+p���܍���n[��$?N��|�&�!fn׎��gy�S��
��m
�w@m���ۘ�g�o����Q���ߥcžV�KZϮl�E~ ���6�8q�CL��o{b$%E����`	E���l�&&������B���zӓB��X2�89>�C��b=T){Ca���vZ��g�y��a�!'�j����)�ɖD��:�ji�r�����9J�ON]6�����8�B��mR�`�~B�8YX"�.����h�Y��P��ڝ�`����rQn:`���� F�6���c�.�Ǣ ����C�ڵ�����G�JG7��e���i.7��;�l���W��g��j�d��+�t��)���/��Ӱ�*f���V�9t�׋�?�o���$��2�|�=Tc��,�xI�].�+���Ao���y�.~���hW�n�l-��B���8O�4�S<��[W1<�4��i�}����N��7r��f�����=��W\>W�Q�l +*z���О<������X�)K��;3�h�yG�re$?+	��%Y�e��4����@H'�m���o����	l᪼�����M�Ñ��4Nj�?0ps�? �;�C��9g�R��C�Ǔ�1�
��~c��
9��}�G��0��~vՎ7�������K��Δ�&�uS�ƅ_�pza�.��s�a���L ��Ｓ[Ɔ1[zG�U_�QB�1g�3m����F��#�ĔQ[�2�P.~Z����+>T|� 0" O:晀�,řh'�t�b9_]ó�q$[}�#u"��6��h�����kx
b�z�D�3T9u��G���r �����n���������h]NAE�����8#���wxW�pN�q��.My7��
`h�%�x�ϔ.t��y]���=��ַ��5&`&{=٥��ڒ1�w����Ũ��X��N��F�,�߷��샠�&�~/��$��������ǹ�:��h?�B�	a�!B��9�G�ć���q�b��ـ����?��b�8b�lpÃF��9��H��i��|U�q��s�%�i{�9���vqZ��/�$[�G�%���#�>:��IT�>w��rM[�8�{(K�9Q��. ��A�7>�����t�Ed|@̜؄y���nâj�!��� �ͣ��Ia�U�Y�;�h�)l�_ٜ�9�߻�B���#!.7	����Zo��&g��l��)P�=�(j5�f�i7��g�ԓN��qdFƷ)����,�,��[��d4���Ni�l�;�e��GX�����4Հ0��y�2��q�)�������n�SC	�v��0^���{�pѲ��n�@�u�`4m�Xe�x0z���*����E���C~����b��k�5 ق�o.�R&l�[[�����ޫ*12z{�1�z�:�/� �W�߂���N��X��������+=���kD�K}ذ�,��i����w�EO!�m�*�L\�N5Bk�Z\�,����~W�$ڹ��`q�$�UF:�eW��^���r�������v2��5�"�*�/�yrm����l<H^��[��qM��v�e9��\,�b`[����dӔ�������v��o�@Zi�{�6��|���\�R�v�ש��|\����Y����[���pXP�LE4�����k%"2�1�L+��m�0���ލp
u�^�𦱷�:��Q��$��$�#�����L�g��#�F�w��r�c2VAXcɚ�7�"}�'8��<����,��m��'�~�^��n��=�ݖ�ǀ�.����T�`DO�3Մ����b6�酠�0���E�����#p��O��:w�҂�otތ�
����D��o�A"��4g澘u�p�v��A�x�Cd".���<��6l���Yu����ě��3�����=����<��:zANn���Ҽ���zm���	��3�&1Z��-C*j�9dvЪM@��{����d�"���"NV�U���j�L*}5C�(H$V�V����!EM����\��Jܡ���^�{�&�E����ɪ���پ��ٓ-h@�Q=�:-ť-�f�N�����w«o.�M .�}@}.��bp�I���hs�q����}0.YPV�ݻ1j#!���-����|�3{۷���A��i�N����ML���L�sר�^�:[��Q0J�`z�>�������_���v��pEo磥d��Q�9�Ź��IG0�sfX�����Vɚ�t����ߕN���"���:�}�%s'�w�Z��M�8�v0
8o$��8Av	��sq�Ɛ� �U��2�Y�ι�"�	rO�?�$N|n�ۃ[�F����$A�y�/����_Pw3�JR ��<@p��ꁕ9*)��U�p�m���(��N�=/�ꏸ(�� ��&P�hL�Vy�:֮NvMĪ�^�42�_Ң�X9
v�Ę�B~���}�ٰ�F	��S5 K�)c�ܓ�89ҽHi�ɮ�,@SO���[2���8�$��C��e��{�' ~V���O	IH��C`Qd�)�Nޯ���	���B[�����L��
����AJ��]	�r�nz����2�s��]����Zʹ�U�慎�|�
#��Y�6�>f��p�����QU�W�-
hn���~�V��%�&L�߀K�j�S�4 't&���iki?� �$�$x�fcI��Y��|O�{���> �/p���<Q��	 w�kL�������H�vx8���I��@�ˌټ
����䖸�7'l���΃��{�Щ�Bhc|���1@E�+#HB$!�%GQ�� ���џkVt
�pH�Nw-�E;���z}�f���c���\��߲��)���q�"^��bM1��)�Pk���{���߆��	�Z��`���ݿ�M@ ׺6��{7�d�ݥ�,�$.Z,Η���#H��d_��f���6����N�p"ņ1��p~��6L��F���0 ��~�"�N!5jYA��J���V�$*&���Q�u�Px�G�3�ˡ�ze>Mz^�n���4Lm�y���w��>�7��^b�Co�Sbq�
��0����B���^�Ò�5�bdu�!�ջy>�Q2�@Ll.��`;�����+�y{%ђzn��*ꓹ�Ќ�c�+Pw�;�����Y^��������4)%�5�1���K���������Y5�0��h`(~��v� ��$�����p�۠��e���/@�gVAD�d�7^T�X��_����&�_�����F�C:C��³f�^mf�r�0L���{e���EXPmk�:m�Ϝ�t�{�&���2H���d̑��Z�6ƅ�T�>c�l�b��.`j����+#� |o�sL�Y��w�z*6���ۭ0��J�z�ī#�ʏʣ�>%⦯h���Yk�x�}pm�p������@�S� %��Ke��x���|OV0X�+�b�aQD$b�u�� w��k|����A
�"/�U�4�Bǩ��G熯��փ+���"BЯ=q��m�b��g$���5Eg6.��T H6<xx����Pg��b�dK`N/��	�w<n�U���#�nH�ȺQ�={Jl�������y����+��� إ��+��ڙ༪��M �6�+,4�Ŋ]aNe�$�#�N1j<f�Y�E�
�N�����(`��aB��Y��+��Fyp P̈�'ͭ��2�h��4r3�!��xh��Wۈ�H����7̙x`�q�2�3�`��a�ȟ?B�L�9�0�nm�4�6TyKT���`�ul@)���iUJ��,>Bd̏��E��T�L,���p	�2�;�N��s$���Y"J�0���T
�.��zW�D
P��^2�����_6\zfm�S�]�B��U@҃���|qR'���'�)�J�mP�kҺ����%O7t���wT�:㚄��E���kO��z�x3˖mf�
�T-�f�����e#�ԯ��C����+�y���c�X�Ž���(]Ih��61�y���w`+="�������A�R�<�&
�d�ڷh��8��R��TG3��p�ˆF�rS���۲/=�٦
C�e��ª�%��B��� ���F�r}MH�| �׾����+��n�ҽ�
�[�i�D4F(�:�!�����I�3�4��]j�a�SlO����ɸ�5�[z[��`�CZ�����s��ʪ���%(�
\���A�Р?���Ę<����P�s:�!{1ro9�ik��%,��nt≤���q�i��h�e�3&�SsWॊ{t��K=u0ub��pf���mM�����0���Y�D��`�w%<�u
�]�A����*�3F��"�t �BTY�I�$62���6�>�F��4���v(3�MIg����@��J��4 �H~/͇.ؒ(�V`g�F��\�FC]B��xv���$9�������:)az��&���`�e�r��#�3�g�s��0E`C��f.���� hC޴�Gto���4�Y�B�-G�c���B�z�#��E�����Y"�W4�������/
�<��/Y���c�AIګ��j�׬752�a�L:�B�f�N(Y�1G{1|cI�>��f�h��V�MB.+�i�]�B�k���٩H
�A3Jl�H ������W�
5T{E�z��X%U����5N�6v̒�?�������H�ގ���2��<x����##BX����+[��ʘ��pj�Q��~vk\�9�}�@��m�j�b�#H>EK�̀e���R��>G�z/�f��	"R�I�M��V��/����A���b��LEx8OU���ɴP���
���=Y#�Ϭ{�n֜�j�$2t��&�?Q���vK=�ܯ��fs`��'X���^]���c/dV�J뷒%6�8�ġpP��E2VˢJ;��]�@Z�0A��
��w��m�� ��z��}w1�A�s��F :�#���PY�3�O�O\�'��~�r�n�Es��d~A�ᵄ�
	~!3�eݻ�s�@ք�>��KMh`si c�F٨?.������b� �3XS�֬~0h0��6s?u�%V�����ɬ�S�� ��
��K��Z�5ЧL^���bz[�b�2{A9Y��d�t`�A�xW��n��wDfA��H%�����7��R����% ��|�b�M����W�
��j��,��SӸ��e���s�*ֶ�� �"+��2�� =	+Wb*�����>��cY�uf�,s�׊
B��޲E��R ��n��R�76>��+���Za�.;���Xk�/���G�}e��kB_�͑�k¡�����V���1����{���H�j��w�2ȇO��6�2����Xj����_\��)Mc5��"q��ol	���g���W�ib��85(�Z�x�W�Vbv$��T�q�o�W_�v���|$��q��[n�:1����%���T���qޛ���uJ�;�Ѯ^"6�Y><�7�Xo��%�
c�������MP�����5W�K���?��@��E�MyɇS��25?�^�{��(ܜ,^���D	DTx�	���4�6���!��E�b�:�F��Hº֦"e���T-5�©�!}< �<�+���v��T�����@��[�f�8V\��n�c�:k����?����%Xyw��r����>��;����k�Mr?Bj������w�d���D�����7t�7prs�^a�d׉4֎Uq����o�gd�%[����`�6�H��SV���R^����ȘA��[��]�R�!Rە�Ʋ�ޝ&�-:�8n��N�S0����P=�QO��(�+��\�Tv*d�K�,ދ4�2�A�iv'��1Z��U
	\!ׁS*�wcU�\Ǹ�W�>^�*C�}c9�n��v���6��ˁ�(�C�p֩<��U��n������Sse:�ѻ�t��v������m
 �����_.Y>>1��R���<T���7�8�k2�]�akc_��a�j���[�MQ�?����f����r�l���^@�����¬��F��DTz�"������%D.����>bU�w_(5���e����u>�|	#�[�h�;�o.�×��f��c�H�����\����Ώ��]��5�eV�Do�MZݧ㾈��(�PTv/d���`}K���ΗO�5�\9����a\���B�
Ê�>R�C�H�ƈrR����}��p��%�ϧ�v3lJQSZZ�f������=AòM#�h���Y��Һ#3bV��X�M��2߿Ǚ�<I���n�4��E} -��o�n�_%co��
j�yL4������8蔕�hG���kn���a��Pr�q��z�i�`��(ˉeั��63y�M����]�	����׳�y�µH�d̗֓G+@y��Ѻ?U�^}�l����w+��(/�����H&��7Pa���u��OO3��Q�*������M�%D����r��L�=�~d�?p��/'(���C�7��`?�3�Pɮ@8�?yW�u��]��	wB��B��,LhK.-�/�~MJ��C3�4x���>��L�&���.n�1�����Z�� K���rGs�ۂ�r(lrSQ|��`�@�VDmh�*���sl��sБ�Bd�g�����T��j�?�"���&?�<���z��cV��m|�+t���5�C{�CQ�8z ����MH H׷vO{�fD�* -�X��:q�<�H��ϱ`��p�&1ћ��*�m�-��v\];x�E�Eޢ�F!��[�)qE,�xc�2ň����N�բ������/'��>~�9�AU�'ex��	�c������ݛ��~�JXNb�v�w��Q6�?���I�\⁛�hq%DH�G�Ɔ�	��$�M���'���.%��C�bx�*�5�zPH��^%rNR��Yoo���6��µ��x5:�� ��e�>��s�.�`qO�>b�A{S��\�	�j���G�T�#�,��L��/��;�|t3jh�(�G���2���C�)�H�k�4@M�*��H��@9N����v�5�M":c3i|�r�yp�`@�>�R/����ȿo�܀��0�� �npS�j�=,�S����9�K�|�]+�Sn���� x�,�~p؅!V�2і��D�]�t/<�Ϛ�.��K�������;�,5�uԜ��J���~�������qm,{�6bO���k7��,�! #���~��St��U��U9�Xf\�V$��܎�#qp7�e�D�-��y�Q���^oߴBQ�:(C?��Z�q`�@n!v"�"nYׇ�`�M��R��)�\�b�|#��ڰ1B�C2m"B�u�n?��sJ�+ߚX�w���.����"$h�fx�R�G��nS)���W?eM�Z���S��c��D~��˓4��j�.[E�����%����>�f�"s{
d>Kbr��Mj�#�z���Q̪v`�ɋ�}�W���Ϛn�����K�G�8c����l��b��Ze��[� S!��Lu�& AVc��QV�NT���tm+v�}�~sm����Ht���b�,g��`9:����������M�gb�����Q��ꀛ�pL�����B�&�3Q��;���9����"�`5>�\��E�������F�_�s��F�"s���&���ݚ�M�
(*�	�Q!Ԏ:���Zy0��A���7�T���6�+X� �AN��*�4c�1���V���V>:\���j������a��}�%'p�_U�im�]0�ݚ/=P��fحh�a^r���|	K��B�����&zѪC_�Zw\t��V�����R��'�M:��&�����o��[M�L�MnO8[m_��ߜh��)\ۃ�X�#�X���#h�@�]C��զ�Y��usЌ���>6>�����O���3(���G�&�pR��:��`�����3�n3�W�z�g���w�A�7�����a/Ĕ�+]��15�&d^#)�d����G:��	'�.:�O;�6 H9��\�QKnON��CvW��ڳ����F��FjWU<�o���	ˏĀ����MJ�+�!�0kL��;V�l�Xt�{��
�J�M��#���z�M��Hl*Q��Q-���Y*��������{ڕ"*8�I�(���%pڙ
"���FP-���c��ՉI��v�bI���t�OH0jDW8���0����Ӷ!S\���� ���XL�	H�/�3�������'z�_=7��h6Y^��x�l�d�T���&�;�%�=V��D��z�/�E�����}i�Ӷ�d��~�nb���ʟʢ;��Pn�86R��w(�c>-���[�F��\m���,�'�*CW��z5(۬�i'�R�<k!x�	cFW��L��d�6���x���J�9 ��ӑ�SP3%���� �@�G���_78�'�py��u7E����� 9n���җ�0mٝ���jy��ZR�=`�JAz,'oz����Wӳ���-Ho7@U�5��P� ����
�$
-�E'P� t+jp}o��rj95+��J�|3.��ّA�)z&��6*�	A��b�1dO�v
N�������\$}�t\��A\���lb>���C����v��(�b�H�e2(ں�+�}=+'���i��U]��㺦$U'�^uÚ�� �^�ЊK�(���.��Cu�ZV�w? �(+�Zu�ę Q�	M��:ܣ/��?<���#�ڹ-��A�����d�A��Vɖj�k!��s���nW*}��X��cVt~��Lb����C�	�X�m�Z���W�]�w,oCϯ�Ǜ��>)��J��U�iwV�S�.�$׮5I�����K �BU�'��2��#2��Ѭ�I��?�[b}��r�-���d�UsT_["G�h�U���֡�f��ɗG���V۰E2��U�n�dA�N���N��-`�5۵lz!iw
�q�g�gP1�W���
 X/�U����anFc�W�J���D3��a�E��eJМ�x����bF�����?Ϝ��`�!��Ȗ����z\�����CQh�����1���m�<!�]AW�k� "/��h5�Sx#�1�,��rP�"��V-���I�m�E5�|��,h�3+]�W��]��@��9����`1Q��u@Žgp?UV�w�6�zˤ�r�ۚgF;L:��:*u	9!����9#�Č�5��b�v���Ѿh�s{�r^�LHzm��;x�M�r�� ({�x.xr�rn~/�l[P��
�5t�A��?���Q7L����R���jC���ϡXU�y@�`I��̕�Yp�o���kj�9����{�,�N-7y��\�c~�^��� =�UH6+���9i[�������`�vl/�z��\��>Vi�h?*����8�� �9�P=�3�PXԈ-|An��ۢ�������k��L��*� $�)5� ����L
$ϼ�Tg�����@oTSS�G��K��28�1��֋����X@�@Zn8�*���.X�:5�&^D���Uן輛�qy`������	�g��~n.V|k��C���D�sl`ۊ��5 ������^�\v�6�����K���ۼ��ێ��+��iq��I.MTB����u��O���H-��+�콿1���<aED�g��¦��U�\f8�W�Nb/�E�
C�ĳ��>�Mݣ�(�,�i-�OQ��w����u��$�>Q����FN�XlAě"��GP�mTʂ%��,xᰦ�|�{�}�q<�Ű�i%�<�`����F�R����Q�gف�*L��WUiF��ff��i�_!dSo�+Lt�$���U JJ��lǑH��Y/�T8�f4f��uyC�����~i�Q����N�9�7"��w+���t�Y���;.�૱ɷ����>��䚨F6��5�Vϒ�Q�=v����gV��2�zC����AOt�L���c���z���ij����N���&!����iV��2|�G	��d;���?m,(�	W2��i��;Ա1UN�X�Ӫ6��:��:���?�6q\d�F��/�`T:�v�y2;%Z�ƌ=J��ܞȺ+��|�F`|3&�i��TqZS}�w�j0hՀEwբ&�'=��{�Q����%�^��p��t����I�H�e5T���1B2M����$5�5?t�F�r����FJ��v�h��'��DO>J��A9r���K|�j��v*��ֲ�3���}G����ͯ��tO�]�6� �sgN�H> ��C.P��W֤7b�I��>4�7�X�W�<3�h��5�W�F��5����F��&����m����aW	�[Ԏq罭��@���7>˹{oƜ��լ�&����+�Pv!�����; h���yO�(��d)�����Q`*FlP|�y��4E��}�f�K�\�q1ɛ��Ks9�� #:vmU���J������[�1�Cߙ������&���;�4@�� /C���jk�Bo� k	+&�s���a�G�6g�jޱ�¼@�� m1�dr	�f��.����#6�<HY �F~���Oz��-Y��(�nM�Ę��e�V���7Kj&E����H�Yg)5Dз�<緢�W�j��m� &KH s��D�_���=Y�T�84�@��^��5�9qb}��������ݴ8k] ��!�:2��q��oU�F��L�~L�tC��a)}�K 뚋�4�<�&�H�K�o�2ZK�O��SX�,�,��f�G�O�*�sN{��E�.܋~[���"u��Հ㲾x�po7�����vm�j�t��t���^tD(Eg�[��n���$>���
u��>I3*-�T��	���s7̖�t|��B�S�d��	#f<������?���g &:be�G}��㘚��ڈ��q1-�`l'����op�l���µ]�Uf���GX1q#��N�E�DI���.Ah�۫-��O$�"ޠf���!��趾dڭ	U��mGd�%!�-�
(g�$g �T�.�I9�Wǭ�[-�~��4v��_ޭ6w>�{�\��l�rq�-\U����fcz�y����G��G��bK����||�d`�:��"�?��%Ar��Fw9�v�0EZ��i�E��UWJ�S��?�|��o#��+�2U��l)�l�����
�h�4'Gr��<4� V���9=p:E��1��]ֈ��S�m��/~	g����/9S�m��Ǘ��j�*�$�ử,��F�=n��J�N���n�:NT�1��,u���"V�5Jāc�_	� �L���b���a`���3�:�Ĉ��XB~"�@�j��4�Yк���	`}�F$� p 	,B�/q�˚W1M>���.���NS!m�<m�7�������%��/l��X�:3=,��i�K��(��X��;o05�+.�慒2���bafҨ��)o��l~�d���b~909Ʀ���DtO�N��E��H7�Q%�	G��I.�3�v���*��sкi�O��}���l��D(qX�=�����Ni�չ�3�k輸�-fR����D,C��$�]�����.�����!^%c�1M�mZ�Z���>�+��'Ǳ�*�ؽ����@��1��?L׏r����������IP���\@CP%1�H�"�Z�iц���u���vhk�Z�2d#����
�8�����%A8��|{���=:� ��T���P��V�"�΢���W	[�^�g�Va��̡|�ڃ����-$f�Z��@�w9��0����natK�]�
�ՒZ|��4�/���QH<�k��4r\�����NǁQ�$�n#\����ژ�[��ɻD�.݆�lVvT}J kX�E����4�$p������)ﵗ
������`�&UD�scx�����������tA��
�K� �|�C3�^�B�
M�;|�XŶ�L������o�����A��+[�6Cvyu���[v;�aֳr�
$�f�O�=�O��X��G��@p�����)\׏�+�nһ��c���q?*�9�lj���[���&z+p��wT���H&�1i���dʀ��Y�j�
+��`�<�D쭸�dN���'A���ӧM��?�������672*�RN:_;<UNҥ)(�[���ݹ�w�i��w��ɭ�66��H�(� E��<#�Ap�Ծ@�$}b& G�53��s��� ��&_��&0?�S�y�`���x�>����>ǋW��G�C U}���G�ɨ��atּ�.u>o�퐗�����AM%�M3x½�����"ߍ�g�����X�y��!�S��$��퀉@�V�`��
���d��=y2�����q�Y[y9�[��iKc�DolJ�)}��eh�.��~�R��+s��X<�|4��OM}��������@��"<�/H�ܨ]B�Yb�y�z_�2��U1e���8�#(y�/LtP��
�4��ʑ�QTj�����J��~F�ͻu7�$��UW�/ƻ�>\eK+X��(��0h+j$u���@��|AG[?��z/x���݋�߹~�������)0NV��J��E�b4ۜ�ɔf�,�����f� 9P��?�2�Vi_�XG='�}F8!���V�3���j'":�_z�5�-�� #�|�]7���fa���ܷuS�窾Pć�oH���94�'��$?�����D'q��#fڹ㛭׼�w����W�}�����2����I��䤵Q����Ս*�5�^`��u���졩8��D�}�S8^��}L*sN��N��=<������޹�׸$z9����X|{1~<j����b�j�tH��"�C�0��̴d{�F�r�/��I��/���1g\Ϣ;���z+�������&|�K�e񬪓�����5�s�'�;�Z�ٹv˷���OWi�d�tN��D��x~�$��F�~�>�2R;S����eϦl�L(��I��A�����V�{�)��	Lr����VS4q�Cc.K�a�� ���g�7ܡ��TR^Z��,j_��R{�8�k�ǽK��R2�*2�J{V��e��+�P(q�zD�������;ZM������_]��J���>절-a@.�b
�����r�+�Àr����*aBn~5�7�|�c���^��<>
�Z��D�&j|H8*�W�O��2�_(e�q���螑�)DAP�������5:�m�J���b�qs�s�ڸ݅�kDfӸghN�-:��9�A��"�x�u����ᑐ��Z�!�G*���� i���2BX����m��'.����\-�c�"���Ҏ䘚���n��U���a��s{�lܝQ���!��i�i���6j���������WC?@7���8]$��?���D���]����9�Y4_@ؒ��O��2�h�҈b�$%���N�|}U��!�C&�1����q1l�v�{n��s���#Cb3,��W�+n���o������|��tg���;�k�0�2n˘U�>��.Aiސ{��kLqw�v���������z���%%a�:K�5~4>����NC���B��L�g�CK\k�5h�g݈`��C.������5�'�&�X�L�`�=�P1i���e)vQފ*��q�}}j��%EO�%x�:�P�b�\�L�"Qn����7wrʓ��R���	0E����kr1����VEQ{A:P�k��bj
F�ؤ�;aFl�2��Ŀ��O���ٚ�*��;qs�� T�۰�
���˛�wg�$-/�aҜ~qW�W:���T��!<A"Aw��8l��]����`�¿��PN�9	��}�ƹ�`�����ٺk21 �l�D�J�vq�*UZ`����͑�tR��[~hБ
�Ǻ%Ex�}Y��n�8����0Α���&n����8[�׼*;K��E ��|��t;�[��O#d	*o�龝 �u�p��!Ԁ2�!��ni� �\�˒�(�A"[�8��l5'��b�OÍ/�ѿ��*�<pg���>- �)�X��=�#��
@c8��mmh u�\>�[�K6(��.�+1�zϟ��jQ��Eኚ�!U�4r6��5�R�#�o�x�Ԓ��Ƥ �<�e�_Al48��	������i���hbAs�C�Q���*�It��7���ll�#��2�����>.����*�����=���m�+_�B;G�\�V1Ż2�@W9b����� 6�(�S�
3Z�|�rwB�ѣ�T�����^8�,�Z�h��jD�j70Y�s���a��Ζ!:,y�=Ik(w�X��'W�m �'�_�c�VjQt�9�/�H��E����C٠Aʖ"޻P`�N�G`7����0�s��Q>��	�b6�Q�]�7��D�=4�0�zhp��T���X�Ę������i!B���zt3�u #��yԖ*�	�����ȵ;*i|v�Q��H��\������Ck�%)d��2C8���:;:Ԝ�L�Ǭ�|5�u���Q���Bl7���X���]w�끕Cz�wW�~�-�7��\ۨC�+����qG��v}#@�1}ưjEG�ti1���+�:�X���b\[�8*?�ܤ�mn�o�9�N��NW�f3��eZ��X��s��\7�rD���o�d��O7��kщ�"���\��X��n�)ZoR���W�N=e��%ӄ����5��ݤū�WP�x���2�������Xga֧�����sd�N��*ؒ�E�~���.���;�W2x,����	j��M��w{����a�T4	�F�Dr��tz������Q�̎��cW�=��uŐ�qY/�?�$(�&`3qDnM"�]��k�w{r�N���	d�W��C6j�/�K�l�M�qπ�mC��h3��̏|�W���� ���NUw�#ŵ2��Z��9������Q͇\���f�jB%ʳ���GF{����?����R���tE��F�uL��!$-j���(\]�Er ��J<P����E/4��΋�X�7�!��6�<.��+~��q�1A�<��l0N�4HND�6eM�a̲��q��xhW�}����3�����zy�g-�iᑭQ�}��ZP}�6/8>/`�����c���V�Ѐiʪ�*zڽ?��!5�MK ���r:�*�`RQ>[y�
���f}�Ϡ󱏇�Z{�0�����B<��~+�$�$-�����=0��U���*����^��48	;ܸp�p,�/s^"e�QVE�8������`�a�@��������hJ(W	�%)!�4A�`�2�"��X�R�R��'}���K����]�0�s����}r�iW�����km�Y��'䉒VQ�R���ͭ�2�y�\�3+�2��3��GpM��-�$[�l�j>c�olO����#��$;60ܼdg�ʸ�#|��
n(�j%Ĵ�1K�B��[ �ky�Z��^�D�E�J��\ru��N�e��}�;8�p�`��R�)��S�~��׌U�H��`�|�p`L?C��~ݷ�����$#����"=-���Ѯ�WgS+{���=���'�
sA�:�Uap���^lz�
F��7,W�5*��/���]X�>N�˺j)h��N/�.���`3;��X}�v���1ۊ?�s��!����l3�b�K9�$�㹵ފ�����i}���C`�6[d!Y�ۈ��������K#�ކ��S�`"�Ĩ�f�~�I��s91l�f�yGxH�C���K��<��A���
�[H��R8WL�/�ڲ�ǆ�Vb|W,B%t� �c�_��Ѷ|WM�
?��)���Hp�)�=���hD%	�F(mk�̫��J%������������s��B)OR*|lr�n��X��)�g��.��D����te�2N/*�G��j^9u'�����'5GB\3+��r����ZU~�Qb�Mݟr�R���9�s�k�5�=��V�Z�x\8v�h�1X��4��>xrBݖD\纩5g�̄u�ZnZ	�uy���At��|Z_(�^�;���&��Ȑ2Z^��������$�Et�iC[ߙ>��²Қ��ĝԐ�}'ѷT^�����< �5=�c��J�a蓰�B��c������>��r��}dh<M�O{��O\ᣝ�T-hy�NRC�#v �e&Xmw��N4&Ս�0�F��e Y�X�+�癒݄�$�����EX��>���IH*n���v��Z�`:���.{R�.��.�;�����y�h�/d?Ū]�ʁg�_��V��Bp'�@�q�RL��3�"�������&�.:�E�D�	��%D���}mt?�F��B�ZY2o��).�ѥ?���}���+M�An�]	�s&k�!��	ثM���K� ����B��1��nx��@З�X�J)R��2­N�Z�@�R�2�et�x;Q���d�S�)��`!A/��? �Q��-��3:>�hU�c�,hS�^���j�LJJ<�e����?�H���WU\=7��Amf����ܐ𴦯��h�fъ�s�G!�+����3��� �j�H�G���Ū�刮�Y7����g�����L��-��2�6?�Y*���r��6��;�U3e�MT=��u*F�0�GJ�n��MP "���[8=�c�'�S���S��n��t��j��3GRv|�X�)�6K�L#���Ϫ�&�ژ�R��ҟ��mÅ:�� ~����\�d{��H������K�'
$ݗ{��G)Y�({��Re;���s�~�� �T���r!��_#���;�/{�;�����ruig�`uЀx�g])D�:��1���K�-*eQ亠 _&mW(��f$���H����h�����eP0�I���>}�7�ٷ�Q�V�[V�ɼ�d�ҍ"��=0а �AN�������s��n�]���n�6��ƅ�T�m�7�C���uS"p�=�~o?'M1����r3��u� $�Y����bH}F��}MkNv��<�rݧ����ƒ��͊ۥo�b��풾&c��4� }��&��&%��b"�0��ʪ�p�#��U�&����5úM��uQ��.�� <��zm���3_+��N �x����2UQ&ѮI��\(���O����(� �ڌ�钬�{� ڂ�E8�ߍerP�c�<��q�)���6��������<�O�W��R��y4��?�۽�[UQfN����AuNY���\��S_?����<�w�>���������uY<Mw����F�^&�L[AB�Ӫ��F;�������ر��uMv��/���Cn���P؏�z���v �� ���B�`Qi7���R��ވ�6�7B�)���ek/����%������ �fqSW.XFی�g_�%n�*r��|����!��V}}=Q�3�5���:�R��C�yb-�wT޶��1�"K�(�����W��/&����<�z�~��ZH��SO8R�UWh�~�E�-�/(���ԉS��Ͽ��<A	(�_�����䍉{1]�W��^^�O�/ P��(�#��Ԅ@��.� 2�ښ꤃�7_ڡ"Ǜ��Q�ZT��6�=�i�S,G����j�����<I�j����D�*�����+��[���	T4��+�n�,n ST��܉ӃF>N�2�_}��6B,��?�C9���l��55�V��'�f_f}!�}�����M�a���^@!���5f���)[����ػ8�Dۻg�ʿ����
�v���[~()P��L!rȆ�vj�6\P�h� w��#	n"���1[g<w{�\�{`�	�x�B c_p r�#���[����8��!���ǭVw��{��O��rY�M������M��~ �vRމI�h0���@��V��͠nu��8p�U%!�e5BP��F��N�eB�\��w��#��0&j+"����;���ɑ��L�7��me"���g��*���X�54u_�ʈ������޳U�^᫩�e�����)�� ��8�j�1)?@���V_$f��0_�Wa���2p��ӝ?TF���[�����n��z���`�-�<��=�r� � F>���P��#��S4��6�;0��Y]�7�xAZ�Sm��մ��w�(	Hd'u@h��!0�h��]�5�?�Ϝ�L�'1O�����J<WX$uԽ�>ƭ�q%Ҝ}�y3��O<��{f�9o�W�>���/>L��jo �o�E��K�u��{����>�;��vԖ�M=�
������փ�Ñu��&Kǃ��ßBIV�����d��c�y"D,�~ݶ��W\��� /Jl}���xFA��C#��jh��!g�j��䛌�P���y�n�#y�5D��:��1�<�Fw�������:բ4W�o2���>t"�i🷥�Q��ygvcP�����$%��R�&I�Oe����)����t��PA�UU�Um��N�m�X�ײ�N�(9�Y�S ,�89�o��y�$��"�D���1
7���9ĂC�B�W�7	aFKP�箲yYTˏ9�Ez��EK~+W#�f��	f���>Φ�C�� ���������7���MZs]�8�~��^[��{�hiGM8�f���ՊQ?7^�Ė�j
�AT���U�ތsw�V}���_�/��4������0�\�w�N�#�>v���Ln^���)�e-u�1\�^���}'P��G�sB���Ӥ�2x�Џr&�j.��FA�aʐ�Xd-��`>� L�y���=���9�a�r�n@�$�FĴC2���}d�C��/ ��n�u"�a�U>o'A��}�a��$2��v�L����_9���ĝ��4���B8ċ�市��[Q��# ��G����No��S~6�%&BH	l�`h(`|��w�JA��J{R�E��2�n<��������:��}v�H�Z��魑��b�W��3��`2��֒���fM=�*k��I�`K�m��H���N��	�)����^x�b:l��>��Y&�b���Wؠ�����kw�j�D����!��	�hV������Ps2�>ꋢSp�z����Zv��Y;�Y!�6��k��\���ʦ���2���2����K�)�:�M�����\ޯ���}�����v��.M�'�����Ò�5'�^ ˒�ƈ�M�*��a�t\o�q?O�/��ʳ��k)�}k��%)/w��t۟���FڒI�yhcl��@����FE�{�7D�*�l�,��r�Y�렦��^gU������q[�L*M���ȕlEK��}� �*F,�������B�`�jT�̗�Pe;��h��t�[Z����m���D�E� ����(�Q;�d��W4���S\|��ܬ ��-�!�3�{'�����~_E>�Y���s.�`L��%�����{<t� l���T���A��{Uf�J�աQ��n��e�%���fЯ/͘�F>�;⪃�.��ת��0L����w.6V�]�/	�p�̏�s�VH�����G����nX>�g��o�C�m{���5zbn����/��M:�X�r[�M�`�v�!UF���I�J�*KuΞ������%q$�u�
H!@f˳����6n���K-s%BR�a�������\y�ݘsKp��{b�[�O��ݗ�� u>��][.��ˈ���Dm3�w����U���*�%��MT&죏�&��-�Fu�,�r/�۪�Io֦W8�#�ת�Mp����r �Vp3��f�_�����^(��`0�.+O�����H��^'nŉ��$:�!K�v�h5rM�Ȝ,�B���weXY�Ou�����b6�~x�;/���e���ـ����q-������f�bt�9������V��� �!���[�������Z�c<�=$�=�C�����\7��oL��*nx`3O�|8���(�\/��d&1
-:B!�Y,��ʘ����o�B�zE|��79"u��9Ly����m8�\{"��[+�:h���u�/�f&���L��Al�f_��������m"RZR�A�c\��E�<]�D�KW{>3�������|����I��h�[<��+.�G�{�6�-s���9�I��d�Bk���w�n� f�Z#�<Zzn~�&V��tI�K�D��Jr��ӳ�"O!��L��?��V�SQ��૏|�����|f�>R�Ť��b���|�H��6p$ "\�پfZ�X�A�[S�X(��r;�y��N���ʏ��f��ɸ��������͏@8���'���&��l4�SSZ;�W���PW��wT�}�!�ɻ�AuB-����+�=GY�b�~ j�D����E�^EҞ���y�>h�3�t�����+h@_;���4�.=�BO�~�w�����(����n��{-���j�K?�P��ׂ���F����-�+7c�Sˈ�v��݅
|�%�w�9(�~� �4�4h�{���Inn�-����-��������{�[�Ǚ�+�����.�����Vb�nӾОSN8⑜ϧG
�(�y%��Í�Wf�7��>��9$*�I!LZP�I�t�a�V���ݪ�(?�Cґk>a��$DAo�֨�	D*���Ĉ)H'F�d?��͡i먖�$�dh ���>��%L��(ON7��(���M
�ԙ��͖�XE��=GV���WC;�W���;n_@�lu�9���K�˼pƎ�S(����!K[�^4���6!�+�����
 �^�L(����E�	��\<�4�-�kO$��qV�){瘁\*GS7{����2�x��2�3
(����Z����Mۮ�"m�^�0��he��쿵��cLB�b�"q�N�r��$�h��*�`��xhh?l�~�f_��&e����L��>Lҕ���n=	�<����=x�������g�9�
�������J==�|K�w��ֳ;�\qD����HY���/!��K�mq6��(�'�_������\�g���V�L�̪3�>��`FYO���w���S�����.쬖驔��}��v�|_IP���}��ď��k�}c`�\jfJ�AR��|m��8l�H��Y-�)4"�-��AiҘ�z��	yYw�G2����/:�"Dݐ-6�K��S�������xb}����m��T��|���:p����yOҪ��M�����������0H<��ܽH)�{�Z� *Q��2
��WN�z�έ��佽����@0�x�6x�6�����X`T�l�Z_@V�,�fYDCB?<��>P!���%���0W����W�H_�[0��-*ȭ,�+��'���<��}%Y�U��3��҆Pi{bV,�����p�y�H�
��V��k��]�bޛs+[s�^�n����o�����X�\��׽�
�B_��~��Zv��?gpg6� �l,�}~�O�����G��:�h�_�N�؈M�	�S3��N[?�lb�w�M�և[�%���Y`����{?�%�hz��)�n�Ƌ��T���kw�xn�P!X�Qt9 u��!�D�� 8'~2�C�3�A��Y�;��w��C�`��,|�javp��<���/�u�h>�ʑ���c����%Nl��}����Ԩ�xv�ʩ�&���o�~��xf��K:�W�[����ί��cq��yk���+�T���u"�Kac\�_g%4�D��Q�=�IA��m��A>2Ai5���ݒ�c޼Q�<�� ��-�TM����A�nV�(�r���}�ƛH��_>��t�kwR��R��' `�u�WPw�c�IIv$�&}��ѥ|[<͘��lPtc˫:sm��B�^p~��5�@�o�>����XI-L-���=�!��ԝւy�va�V�tV1;qع`�Y��w0��r��9�=��s��$�u�l�UƸ���,	�QC�\�~NbS�^9�:~�*?j��W�F,[r[�G@���KY4odS"��O�s��:�;�����F��z&z�<�#Ч����	���X���*7�5�k� �Eˤ�G-�9OO�Sv
@FS���y�����E�հ�;�D%�����`��T���Ng���(�35ix`�J����(6���6%����fW9�<b��h,
p���u~�P�ّ���N��A�v�lϒ�9�O	[/nN�3��G�"�X���M&���Cvw���y��B��!x��Z/B���ب������n_`!.>٫F�UG�|����v:�D�mc�=2�
�&���z�2��� �D�U^R��XW�lB�ˉ�;�Lsز�s�����M��v�Rx��Z؇~��ڎ��LسȪ[@h�f�*i8��Gm�=<]C�����q?a�g��)cR|��/
���d�-�xM�B/?a�qS����?��z����Pt�.B3Z�#w��-��)#9��<·}�i��C�(k�>�����D���A�:b�-sqjF_$��(JWDv=J�w"d�߬U�1��dڸ����0����m���j��|�%���hG1����{�?���F�9Oє��0�Nkt��F`���jj�z���{���'b	t��Sg{轥��d�}���h������G:�]�Я������#����q�̹��%�POj������^0-�H.��c��_�g�A��Օ5�e�}��%���FX��)c{L���>w/��1���ɛT�����5�%U����ܕ�N���@ ��*w��o�}	l�i
��'��n��c�p;��C0�rYW�qm� �W@��ʎD����X�>?O����w�W���"���,Y}�(��B���{;�ʘ �� 5p[rjl-��W�=N�Y� �\�.�e�U���A�֯Tp�}_:>�#�NC�@ ���5Y܎Ś��u�zֻM�t�	�z�k��yZ�0[����X�B���L�/A�, ,�6t1���UuÕ������x���{���eCݎ��ר��P��uc^�ލ�d�RLպl�8ģZ���B��_rB�ձ',@V�����7[hF�7��鶏�;x���nE'+��P֖�4	4z��g�KW�\�p���2�1~�]��|D[>��������i���F��6T]V�N�M��x
�t"~*��sU{�~;�PD�$�`Sa����4$���#e�żK8�
��K�F���t�>���y�|����c���Ew�.��:� k�I�������ƅ�����>��aX�2�=;�pg�:D���*4rJ@=b�8�Go�u��ɹ�/���5��F-?�as�W����Ϲ�1�y�?q�ƨ�3�l:��Z]�AӲt�N|�̅��'@ؙ��8�G�6;@4{��@��;_Z���^
���ŝ���r���|"��m���0���u��nc%������6�T����qIc�Ok�P�5�d�r��:�#���J�ލ��~��&��SԱ�ގ�(�}�D&� ���u��xʛ�$�
���p� l-����zM����D8��
HG������u�BQ�����լ���6|�x�X�h�����*RLZ����h9,P�*�w<i���c/�H�յ� m����6t�r������M�I�y8�ϙ�����+P^Y�D#4y(A ���u�t�3=r�rb��mu�|�د8�ST�XВ�\�| ��ȑ��@3���#��t���?,5&�n���G�p�ԫ&ÒW.��柨KS��F����"
:ca����8f,q��v)I?	��-=��z���ˢ���]2&�����禔�$1sBڝ��7ѽG���RP�!B�t�����8aݎ�7��(�6�_���2&��Q����A	�.A�?e�n��k���)	��ʻ�$XNB�-�ͅ�5���j
Yہ�c�XH($4z�嚹�;\�7�X �-#����C�uU:�D�镄�[�7������Ϛ�V� ���X�;`��*�P�j�Ԟdc��V��H�P^D���JR�ry�á��
���؟��T���rjeᕝݘ"��w?��緅5+�*�d�Vn�&4��t�2�ǎA����++�Z�z�5�s�Q�v�d���Q�[ȅU��M.Fܙ�lW��L����u�y��̾�PD��Uh�$>���.A���!�}��(�*���l���1�:h�9+�+m$���\�Wc�6,rB�=	�T����E���:��9��ALL�yM���;����f��ANoW�x=<�MHU�-�dj'�^��Zz��7E��KΥ�;ޣ�$1��|s6[�����"��zN��Hp�{�A�l[�;��}�vE��ΐxԖ����U� �AO e��K�-mo��`��;�pFx�y�YQ[��a)�s�{��M�i��Ez��奱�1�6y܉uN���U�?��F��~�JW<���2��o�n:�x�qr�I	q7��c�3WA]�Bu�fZ�Q2Ҷv�������l���s�g�:"B�����.c��w�P��?���f�ɯ	��_.!�ߟ�I��^9�e����o�t�}r8� �^Nk�%:9�ekڙ���9�_�;(��vڟ?Xk�&x�ޣ���a&�E0�gd��h�7
�\=t�E������k�S�k����D��B�`(S��T!�Wg�!�(�}ƒuK޸^��ԟ�|�ƹ�R��?��i~�Q��3S�x�R/�,:<�Éb���M����M _�K�4�ݶ�+1���%*O+�\���e��ľB|���K���Ү�½{���uD*̿��z���L]��5+���uE�Ώ���s�ȼ�b�W͹w�d��/)D��[���J�[>������n@ze�5��#Y/���I��d�`L>�Dy]/M��	�KPg��@�Er�H ���^ԓ-����vAvɳK���qZ��pG�v��5�QpH����>>h+^�E��*:v���Y�{����_!7Ũ�ɵ����sK
��}���l͋��.�u��g��K���OIA����k ��TV��ax�;{db4�+I'�R��L>P>"����l����{&��>FU�"y�������m���L�$�Pϧ�9���<-�'!�J�%����.�x��d)��?RA@��ͥeÕ2ri#�Ѓ&��X�`���NqH�F�F'�̪a��>�o���Tl\5�G�����cz��6fng�i��"(�e�&����݋`r��H:>oc���c���0�UݗE��~~}ߌM���ۭL?"|���*�ͫ6H������.��5 O;�j�9K ��Ao��V�s��ġ/���q� r�~�
���{��ۍ�֗t��Y�,�}'|_�,��!��M{z����|�� �-"��q���p�K��J�&P,A"�N!�&*6/r�K��g�l6H���Oɮ�]\_
BB<ڊ"s�=>	����rP�󏮶��~/5��ɻ��m)�!&蒼Qy�����i���};�4a �=q��n�ڻ�[�U��=R_hE�a�[Q&��+��}�����~�*�7%7����>�R3� �S�ܕz*7��\eX�3=9���n�_�p���z�7�a+���O����8���l�<u��KB��0�j��ZFN/As}��}#�����:oЭ�B8�9����t���Ǵ[M�	�o�+�,T��X��-m��w�q�%�[�5D-i>>�]X��Z9?@��.�o�+Y�Y�`��[+S*�R�Ϋ�ؿ}�$wJ(L�+q���]마�7IG�_�V$��͈E0
Z6�um%4�?`:�XV��(Ӫ�[���7��d�}�w�W�ֈl�69��.Xc
N,s�{��	��m0q�L�U|u�7�g	�����*A�F#�I?-��${G���L�-[X1B5 �� <�s{��f���"���L��%��L=�&��?�2я�GS�3S"�T�9|n'P9Ҭ�W|���P��j7�
(	�aerN��#s)����;<T�4Pg��H��B�v�R��4�W�G�E���PO�:�lrU��E!(!2YJ���B�Ϗ�	)�n;HK��vՆ�S�{;�sҾ���v���7����'�
@��_�bنժ���i�~���m]$�.q�;��%K$�pa��ڤ�������`�W��s3G�ۤ�C&�r�2�����	T���M��4wy$���s`�s��Nx��0���q��7��GN��~����#^�lsX����`@͘H����6�$���7�A|�nқ��q�	�|�� .�*��P����0���QW�>򂩐[}�D�s7�yä���9s)��ή��8��L#��p1)�`L��9Zk,��-�A��E����.3��m(`Fk��F˧������qZ�2su^���gAxk2�+��e�V�Gw���{/�ڼ[r�k^��t]eR;�e�I�Mߪհ�f��Kh!?~�xp*�Me�o��4#G�<ay�S���������7G	�����:������r#����
����}n��!�q���5
�T��c��[Us��o�˿hE��Oê��!h�4���c|@̫+��3�r���)���(f�nG��.z���jRB×!�/ɡ�	(���ab��1�]dI}�.!�C#_�`UP�b+��t�?1�h�tK�lj�'�/�v�����]���+��*ꋘ~���4��"}K�	Fqo�W�o��҇�}��5�#"����'�� ����$��͸����[W}�����B�9��ֺ$�{*�+m4�Itc!Q9����:'��z`m�NAU*.�ʶy���T��\%뭢�?���8�g2�s�:�*P����0tؽ���8�U
/����s}	8�6=S�	C|y��VF���h���2��%J�/	�L�����4��F�MK�o_�I��j��W�o�����4�4"�a�J&U�}�Dߐ@�nc�>Tp��,��A�����u5��T�����$[����A��2�=��ɖ�΢�D~N�����AuVL]�� ��30\I�"����Ur�Y�=96��"���oUÖLػ1'�[d^u��*)�h�+����L���*>c0&2id8��C?�c6�En����	U=�ӫC��4
2��D��(��m���!o���
�%�ہ�($��(�`����܈R�DbGC��ġ�_����GR���_Ҋd�� %Y���H=�y�=ͧ8�/M�;#E	*��P[���D\/�1M\�ߐ��'����rE����F����]GA��M�ԩ*�h��`=H�U���in��OfK��D���hZ��~QBfΖ�,0�D���T����n$�%��| �m�-���^sT|=ge��@G���YI',�,	��G������T8��:��~�b�"��65�5��|�U�fM�#_��E�ǄnJ���$50Κ��kl�2^
�)���j��%�=�,�g�� f�2kTP?u�W �L3�#g卍��J"�~�z�GD�Rc����	�
l�
�a	�~h��}��0�.�������V���)�%/3A8�϶[��������LYF�2W�VkA�`��/d�s����=��W}����
V9��t��'������̆~�J���w�l��	,�7s�a���"�3D��Q�Y/��-:9N��0�8��J�2/:&�p�ge��K��=R���5�9���M�� {�Bx ��éQ3��O|kM� )���:�^�	�;�OP�g�.x��I���޹c_<����3��Ύ�9��d����"p
A�u�)R��������4��A_o�ل�mԌH����:x�wv�ᒋ��?����X����h��X���sb�İ5�/)�4`^�&��!X��O�B��8�b~�d��xv:~��f�R�b�E�H�A�C��� ���m��c�1�d��Q9�u+����حWS��O�Y?y�(�9�˙�(�y�ZO2�.?���h [���J�5���e��5}*�c&f�d;Px���y���vp�]��Yx�N��Xj�J�mV_~t��z>�0�d!�
�9]6P���bn(�'M��{36�Оa��w����B�����~���O:�g�P����w��G�Z�ǖ����M�:&}jǐ�׎�]�Đ(�QQ�� ��tv.t�K���'/~����f�"�a��])ד��M'�J�4�sr%���n��F+bf��L�$���hz�e��r]�ѰEk�v$�.0e��X?�I]���x��Oa��gWE�.Y�/A�6����0EH�!��흑%�
�B�= �oimq�5���ҹ�U�YK&��o6�ӻ�*V����󾜰Kۑ���6Rz5�Z�k��j�(n?TE�������7t ��<���i�'q��Q�v�oir��A�J��j���5���"V�L�׬�y�����*W-g{SH�t�1�� C�9j^k�\>B��'W�DF��2{٦Z6i^TM��2&�T΀d�C��]�6�BC4��������;.|�s�����/Bŕ���+)m8��ΕHVF\��瓇dS[7w��wyPb��zt=�\��G^�.��g�O!;��1;��ׅLBvSf\��{F;��J�5�LHnqL�6pw�7)(8#>�o��9�Up����
|Y��<}�Zf޳B(9��a�zV0��K`8���ڋ���-����8��Q} T���KR?�1D��.�"`Z��~.�H��
�p>�8v���#���b���p����y-P����W+�s��j���"��`�ߥj���F�u_�Wh�\��	�3I����r�,.���NJ]��1�ǅK��|q�3�(���ᩦ��
Q���YW6o�B�?��a�A�Y�L������tc��}Vw��t�r��U�ӑ��H�Nu��%G�>�)���뺈
E����_C�|z6\ɧ�\�՟i1Ղj��.��kRY�+l��޴� 8��A�����J���|a~�қ�e�DY�Zm#��{��_s��y�
�f0��7�!��#�x���ܛO�Y���75��T�W�]�p�K�a:��£'B�t����.��&N~�q^�ـ���Y.�n��6
�0v�ӎ�WU݇�g�	W[�&B@�<����1U0(P0�
��*ŇY��30�˭�|,�]fϘ�/��ӵ[���'x�͸���2��\}$D�]���@�6��]���c��G+�����:vX��<:�������6DlF��qf�7}�(l����o~���ִ�L,��Pz���ːuj������&�H���j�������ۅ���6��]���ER3�o"�ct�
�Mc�2L*���̭���]��t�*QB�yVˏQnzD�|#��j�S�ۢ�L8���_�gx
����A�YGN`����xk��c��?�����Ί�&��V��굙e�<���<�����j�-F�y�(�ׂ���K�N�OFͰk����P/��-���qy5S]?-��|�U��},��bn���=ֳ�>l]+D�2Y���[�%��-C���Ԍز��h�0ȧl��-��+�v2�ͫ̔[�m��݌�K�A���S�J�[�Ԡ�ğ̑�H�P��(
��=�n����?���^|�dԩ�Y�q��~�<�6й�3�0�NS�oN6t8 �>3��]b6���m��e(�(B�~���'Gc�<�4ЗhP�8C��ObGa�NP�c y:����g�RN����)�:@|���o�E�|
�'��#+���C�n�˛#ۆ�X�3��l3г���	�.�d�x�4��2F��q>t��ݳA�S}h�N�������h�w���u���yt���Po� d;U)7"�Q{w٢��g�QUc��8|S�֩b��-�.G�Tc�!2�˚)i�#{S��3{��+���.��R�?>��.7�+�q����1�T!/��ޓp=��=����_^��=��S�"ĸt��
j�6v)Bv�|�´��"N�E^ܨ
���҃*�q�b��1:�b�Ԓs���0RK}}�)�V�ʷ3�_�7$��S��sW��yE��xv�����^���z#l���+��<Xi[�A~C�o�߅a�{iQ���s��HI�9�8��T���Po�ֱa@���$
>ΐ�Z-wW�51��#Hb�O���3�wGܢ@ǯ?/U}pD"�8�wYQʏ����p�@5 ��:t�C?_Z��R'.L	:7�Rg���U4h==�� C�&;��M��<�B�j�;�
���o�	�� ��RÔE�Bb��n>���9Jg��afKD��3�C(p�)i]˫��*�}Q��̻�p�V[�u�-;P��J7)ӣ�*6/�Q��l�+�t��"c�-��~05GvPW<�[R�� �?���ٴ ���A���C�#i���V���n��l$3� b�u�pb�������ZK����lǁ;�w[���ϦL6/�\��pS}�L�78���Ǌ-���V�9�#v�M�YkY݌l$50��h��u�����d��Rj#���~�v���2���!9<$k{����[����S��N����h�1��P����H&Y��6<R4�W��9������ DAȁ�Zu�+o�0�?��nA��F'��\ۯ0��R;ā}��?�vod��𯫊����X#i���"ٳ@;���΋�x���!�J
��_�5�C�J�,��B�'��6 h� �3��cv��(Y�x1��|�����1�kUjbĺ$���*�rſ��� ?���?�"���D��$%�7��~�8��'@�@$����d�TWKXar��S;�>�´:��X�� ��R_��c,=c2�[�0��O;q���3tƁe�3�˴"���2I���>I��%��T{�ݑJ�0ܡ�إx�+�M���O�A�-J���s�.�P�s�u�Q׽�tQY�l�KM�;�܆S;òt��������Ž�R'����`��S��g-xjX::B���<M�m��T��5(�D;�}Ã�WS�,R}d�a?��2�\;س7~��M>V�X�՚`ErX�~?�)j@rh}�����̨D��*.��%:�Yӆ���O�r7�ӿ�\���Ls��re�q_�
6�Fb}��&�=Y�q��F��3��Uj��cY�aAۣ�\��ByÌ9�m�'N�KK�Y+P	`k�d_g�������&��D�p�J���3��lA$��Y�Z���`����z�0�~�1��I��9�7�J]əX54�¦��˲w;����]F���B��J�m�뿅����U�t뮷�}��ܠE7eԈ9Qg�¢I��7n�Pf�q@��X]��;��'��_vЙ�8a�mWՙ�X��!6e�߼����_=����'��b9��D~ �
��U�$���K�/����΂��+���*��cj52(�8�����.�i�st���g�?����#���x���[�r�/��r����w:)���H���wI�cp��%�r�������'��͏ͤAgO-�on��W�g�A���FQl�J��v�	F�d��Ћ3�T�b�I�R:g��]�o# �SZe8��V_��Vn}���ԮrD��IzE+��!�N'��7�&�u0���Q(P2:�ui��b8c*,�]��`r<�L�n{��6SF������
�e�r�G5�*ό�5w�l�h��ngkM��BY|���o���Rƺ��}.c*7�o+1Š��c�$R���8c@��%_�,m��6�ŝ�8؛4�uM�#��;_�zǡ��H��Vnʟ�ƅ�>P���0�'|�9���@��`�w�
�T_m>��e���6�	��m����oAj�tXՊOX)��Dv�oU�=Y&�{,��IKW�ڤ���'Q��n�����~u݈�2���p!16��� ��r�w34vX�~?�ct�+p�$�~4n�9�|��>�B7k0s}D� I��|\�<�����I�ͷN�K���(�/��*�/ԇ1���H���]�R�w�� �&�@q�����s�r�j�>�&ķ���߉K�:��'NX*_J?`Wҷ}�J��t��PWOdc�p�i$ӌ�\���f?E�qtȧ�R��_>�j��]���I��;��}�6��B�6Q��ޜ���m�Mô;�Ng/���]�t?�,�c��+�{Wp_R���~Lh�Sr����A�����3��_��3'����2����]'���ә�/I�����\d�ǟ\r�Э�avz�ڸU��� �
6��RX9[
`�rR�1����/Ƕ�u<Gņ�Q$}�=�ТJ��j�����z��_u���~j����4q��
�2^������;���k�7�-��x�ЏL���8|nte��z 5M�����,��b^���.��y���"�$�)��qu�aT]��C���}�s�X��^�H�$��ǹ4�/\�M�]'�a�=�ƼX��6���K�L`l���by��/T��~k��M�fo����g��JjJ9��X�Z�p�BŢuZ)j��l_^,�ˌK'y�ج��@)���O�㧆=AR�E�f�Ls_�A����I&uM�'O���({�v�@"�pp[y�*�%M�9l2�-�
n�����w����Em,>&�[�lx	bv5�/?ܙ�y������^ ��ri���p>�q��k��e��کP�?n�
�@K�%d�t�6' ύw0Dۻ�ns>���
@U��,�y�Pt�C`����x���9X���+*�Gm�lNZ�V|����^��A��*�ӳ�7��N~
�¡g>����=������/�1���	`�cc�r�Js�;��F��C
Գ��7�ԮV!	E���5��:,Vֻ9���Fz�Rn��{�ߝ�.:!Tl�ۋ�ʯ
I�ǆ�\���C_���+6���Mj6����r/u��>}�y���>�5m��&��/���A�=Y��C}���_�_��p�M�����[���[�C�B��\ۮݹ�|k�����H��ʽ������j��3S�p"^˪x���i3��5U�z"��,�W��&�g���JP"
��~�Ln���t������̊k�YU���CK���.Ǥ��a0���	�q�ףh��Wd6�7�O��ay����ы�C�q<f��̊X�Zb�ᅀú`ӳ�;����I��*l	m�f��~�8��N�sש:`���N��m|��zYHq pHK�Ih�q ��72�.rݹ �t��K��ϼ����Z���2��r.05�5S����p�wf��&'/!t�a1ߠD���CR�R,%�U@Ŋ
�+h��(�vw�P���Sc�큋B�w!z�f�%r��`1�I.�&�y��?������bC靇r��GCLPQi܊b'���q�6s�c�D�r������c����w|��2����vR�wu؋���ZBk�&���o�z#D�O������U9b�A^E�&Ճ����ȧ[P��b�!�s%c�A��Ɍ����%�.�c���X�{iR������(����Tep��m������w�4��{��<�n���>��ŀP(�$��i���-�z	w��RM��z�i#C�[�Sz؎>�E?��w�+��ĩK619��We����Z ϐT�:Ks1�=�����u�^����!��dP	�y_����f�MF�e��V�$Z �n�$%��$��u��F�*Z�l���a��S"dq���N�r"6��j�qY��SĨL�h#����ۺXGa>�<#	s�^�
�EqN@�@�Vo�������!	�HN8�L3'gu�W��͑ߘ��9�������E��ͳ��(��y;(� ł~��h�i$�,-��-���o ���&�`�ʝ��4��$��|.��[�����/��7�=��/���v6�!H�?�9&�S/:���X���U~S�l��Qb���9�RF����G�^��F�0YiC�Y��k�n7� L�f��4�[�6}M�Ck޾=C��T�`{3�����E��[��fu,��,�VHN��O�<�|\���^�1�e8q��;ǥ�eEN���N>{��k���?g��C�"JTq�*:����@R�ূ�m�'�\��\���(���@���Ӊ���5�������𬠡�wE���K	��]��U���̦ Xj���gT��� k�b`=�zB�\S���|���Z�BOQ6ҏ"C�E��(�Y�瓩��R}lh��D�j]E("��7a��fr�k#��B���.S &��1 u厝���T��]}��|!+ް�)�,�A,���a��ڨ�`�1'��&Oמ�8�L���������}GM�q�=i�y@���W�t�i*��Ǩ$W�&��ɶ� R
5����xo-��2�۝�K��X����_���'OE��s�6����Qc��VY��N���Ш"uh�w-�XI'���!?`�{v�i�Q����0dN�,�"�V���+�PV�M�ڼK�jy�`钯�<K�xt5I�|
�!�O1�����L�8���ȧ �k�*� C��m��$@������� \�Ƅ؟!Uk��^W�U��h@Ń�)g�uOl�$���S����h�?;SIr�z��ry��`�%]a:d�;}�]
��U|��)0JU=.�ȼg-{�;U��G{����7�&]Z?���6��0@�fd���Kd� 53�:�%�1ٍ�0c,,bM�*7�Y[g�۷��\��Τ�� N�{�`!s��.T����3�gL�2���1��92}X��L1�0�S�, o�H���.�C�Y:�ށ�	w�"x�RZ� ��p����U����"$/X�Y3���2����;����s�,�x=�:�si|�p�Gʊ*1l�����Ŋ-������1�B�;��G�Ad~�*s�3yR�9��wZx��w���9�G��v�%����7�M+;k��69�#+�Y.d�WMG�#�?�V&P�,���"\q�Y+v�	�J t��%��^o�Y�SBi��=j���X��X���d��1�0��MK���,��fu
��_�gт2�ʰ ��0e���]rz����(���a/��Ե�^��4Vȣ�hU��r"Cv�!���V�էC���5!�A�ѷ��ջ����q��77ި�F�)Dca�
I[r�Ҵm������ �$JB1�WS�0]y�a)�Z�
���K�HRUU�P��=�7�4i�Pkֳa�nsHC*�y��f>�M�:g�ۄ8��aө�=��$��J.}S�F�+�;-�����=�Ց�(�r�M����%�x��x�1�/V�^�~�2�[\I^RGř辶^���ԃ�n�U����@�3eŬ,��P��n�)	�,(*7�{�
� �(�mrw�gҞ"+U�-�I|a{�Cx>���� �$gO����$��P��$(������� ����W8��}�k6�G�w1C�C�/������++�i����6��\���iQ'��oh)�K�2���'<0�	0�.s!�$�1;l\3��^6���V�"�7Y�S�ۛ<rf��#�TS��(��ٻ	��)eA�%����'-[�o��|H�6���uoA�:Qu��-���^����,���JD�a�ɻL�ߍR����Ɉ�w����G�`��	�
���u�i�J�"��aA���/1zU�s��ʟH%� dѣ�c�3�"�G�� ~];yB}��YH�b�h���Л��َ���!v�w/go0P�ҹ��=�1|�ˮ�8�<��R���r`��l����.���}�h��џ��.���s����FӾ��)Q������E������X���� Ch�6���R����R/���3qK`k�^�$�x)���&b�ƓqY9����+�-�8���d�)K�l^�U��Z|��4�1��`r"-'_Qe�A�|�����/oX�P�X���F���G�6��=��h�.�7�;��N�V=^Okŧ�S��:��菧�y\0�7C�YT�gc�dx�=��+�y��l-$���\9Ѹ��Hl!T�=߬�V���K�7��拖�n���{����7�'V7sa�3�,b������ZQ��W�Qp�/�)~>�?3)�Nƶ����L�����.��ƐNK/9�t	_����j�	*�,%���Y���(UWX�1%�xF�+�Ƽe��9���BA�� ��+/�n�mG�jxk�� �YȐ�l#��	,7�~��o+_����z���,�T�bꕖ�6�����˧ۗ����42����|<[��"�2����j���RLwd0G�þ��̥��:��Z�.�\>��c��|)��,o?��Qeq#��o7Y�r�nB��x�.�����D�%�݄�"�2�.a�Ha�h�\�$�-��({Hop���`i�x�Ћ��+�j�>���pRt��Yk�E
�F�VF�+[#��?��xr�6s3�������- �|���Jo���Y��v��d�Z��ݱ`LP���M�<jy@�.���"��v��A��p�,�G#�/a��O�"�Qׂa�ӏ����)X:dΏu:_������6h�9�u�<|�h���`�>��-��q���N��dlD���u�},�X� (>+"��:ǰ�A ��*��#I���|9-��C/��tZ,��RQq ��%^O��D�����U�\G��V� �<��,��L�-�Kk��MӛG��'� �R^�S�K��g� ���B G�^����� ᨘ@�} �M͢q�8swJ�����@���A�e0E��aވ�%�9Np���w+�%�GSц ףh�𔈾��\j`]���ĝ��EX��V\
��������)�m�q7�����#[����KD[������s<_Zm�14��ԃՑ�=�Fh��O]J�w&��B�鋃Rq�_�wku �� ���7���6YC�-�N�5�{�y�7r�̗ �u��O��� �6�/V��f���o�Ǧ1 �JH8eZ���.�s����[��w@�[4���@H�0K��Lp��槱���Ɍ��_n��?[�B;-�<Sl+3�<e�ʏ�1!h�G!�-wc[w��5�2~m����a7��uQ��S��+^���.T/�>N��G���:0�n�B£��I�P���E ����k�೭�XBYCU����V���@'�MI{���hA�����-b~=ո��O�{X��EO.�B
��[0rGFB&k�Bz�c3����P�M��9r�벏�1cҫiC�*�[�Fט�D,�!)�[���^$m7�&������%D`�����J} pڀ3+ݦ�D�����J����*�զ��TA�N++���:�i�>z~x̡K�G�c���DO*�e�00$���NX�N�"Qt�~:�펈A*��ޯ6�üǬY��CP���{cI������k`<���5�(��st�KJ���uȭ��%]����U�}u��NÿUT�4
�7Ҫw	�z�t[&�i��SLdĉ4A�g����T��]>��+��p]�S��`��3��aGܿB����{�K(��I%ݼ�arH��|[�
 ����L�9ۇ��s��]������	�X��2����{��b�呠�ӀZ�G��N5c�4�%�'�d!W��|������2XB/5�&��G�
���iT������!�=���"pZF<0ǋ�_g�r�Mو��5�	�2'-������N����F�lxM�wq@VJ�W9����O&i�.#[�H�@��J>�pN�H�H�8�<��;��F���7��?��,1���DY�#]�E'g���_���d�e�O��gl�㒐�[��Y�a����t�����V�EzX�T,�O*��y�[8i��Ӎ>_� j�|��\S��e�h?U�jP�=�%Z�Z*�VJW��9l�!K~����T�ڑ^68bmf24٬%�P��Vr��g2��p�خF`^Uj�k�>��߀m���ں[Z�8�����֞��~���di��_��v���JK��F�['z��'�ˣ�i�r�^ۥX���E.DW.S�w��!\���:��J�6t�g� ��-	���&���͔:�W+�j�;+$|[��e�І���=�!�b�'���M��;zZ�)?y�7jV��8�6�eKBi�8O�"����6�VY��q�Dc,��Pk�\U�, d�(�A�"��I��_�bcWixR���֭�c��lU����Hbr/�Rc	�̇�K��:��ֱMȵ��Z'˴�yrC{��X�����5ZhJJ�-Y`^U�W�k���t"��+@�oz��C<�20uwk�g�y[ƈ��j� ���QD��o��~B�ք��,�jz�ĔZ�y~�}5H���YyG~�����*�՜��S($�:���j0=^�1\w�%��%}o�4��g�[�j���&P��
�O q����!/�F�EX�@���t�oy׌�^׶��S��ҧ�v�բ
1��/��x��w�K��b���`�#�UU�3V�K9�[wO*7l�p?�MSҝL6G"'< ��$���	��\6��:7�C�\iʗ��1\I��N�ŷs�F�--�[X���Bb�=qm����L�iP(d��h�,��*�|x��o�2��6%��_/A���Z݄v�!��I�>�F$���6]]-��X�~(}�C���VA,�V�z�聴�ϓ��'D�j��_�8pc�$�u�R���2� ,D���q��1=�L�6��Јk!�"�D�Y�Y\K�j?*�uy\�.�rnvD�߳���n�K����Fw7��u�!�J� �����w��x����m���fs�YU��J�͸�AK%��E;���0en�|7L�CF�9vKl�B���$T>��Qz�������d�~lEQC��أ�aN�Z3�g%2H�H��棂#�S&< ����ֺl��f����c���ӷ����|���"�N��ռ���{\��_�D�i+va���/@l�9�k(KLo�Bk�ǟc�`�Y�.��/@�K�|�Z/�F�sY�!�$wӞ+;H١��TbZ�Cq���Rj�ex� x���6�	������{��@i@���j~�E%
1W�=+��.$�:�&V�{-ǲz�U������J:tw��E��S�� 3-r��Ogh��Z�͖��m����| <}������~;�}��c"�M�BF���a�­<��Sf�7/�f��r��&���2�
I'=e���T+�5�=����8񑰆�h�摎���W���R�z��e�R�
��Wߝ�����)6�Bt��j�(�!�	i��Tͳ���?f�uB�~~{z�W��r6�$6"�O�.�!נwໆ"�}�~-��b����f�,m�>��@��^���
J��ē��{�s��<^����H����1fִ�d�s�2����ͅ�W�aq��/LE�yl�nZ6�NKჷ�����dL#/Ȑ�]�#�K.$�!C������t��+a�.S�p�P,����WG[ܺ(U_p����9�Z{�ELfו�p'1<���6J�	E8�%�Os���`>�)�C�!/���8�f�	t* ��&���g�vR�7l�g����lV�c`"3,sw4-C�����V���"��jG���nsC��ʁ��9�4}S���F푩���E�+�CC�p�A��M�2��5���nJ)��KTPNC�GG'l�Ua���@-��S?%_=	aL���ۧ�P�K�Ç(q�x�Q~�0����U�u�*z�[o��Rr�ԺQdQ4�r�2��~j��XQC����7d�<�����ai��W��44:�˹>^NrJ�$�z9�z��8/M�,�WYz����˘���x���fʢ�Ⱦ�ԂZ��>ַ��n����V|��}ρ��%���I �K���~j���kPJd��bn䪳l�����tV��i2Ť��afچ��^�Zї�P�Y�EG�`�C��V!8#��_�������%t�X2)|�C��ʱC��H��t��R��.�O5��gE�6ͫ�en��4H��9�|TA�E	���lMHV��	Ѣ�:�cI*p�;�M"F~�x�y(ZC�OM�v�,� �癭� �7��(<ȶ�h����_�sA8 �]��������$���7���`oBUOџ) ��1�����d�t8I�>� 0s_���� ��*�NX$�ˇo	>(F>Z�I�ن���%(M1�|�G�:�B���Ɂ�����=щ]j���_Q�{D�gf������W/c�Vk	��6)���t�P�vX߭Q���z�w�����"�M�.�N=3�[t��3�/���뱡�g����b9�p켫��2�Z�$Z����p{�O>�0�ߥ �b����:������Q���b|�I4�>RT<7�O��)���� 6�ā��)��t�ػ�w+���k��e��V%�P��=<sHLK�t53j�?on�%�p�4�k����H�*��N�[O�d&2����!5�QYض���C���Gx<k��SPnԈ ��()�X�6_���aX�1P+-PA*��4�3��`Ʒw��D��
�e�bW3o��V�L!;u����+�OL��@����|��e#�듳��v���I�Z<V6�n���#��^ɞGr]��~<�=~rz�I��g櫿>4�d��rH��sӤ�S��I�M]1z�=^"���� ����X8�szs��/p	)��:���{7���� |#힀#�ǉ�� �Ec�e��9��]�p(�у<C<s�0&0��tBt��2*���LCr������^�'��;��Ü!�6��,oU=6�	ē�*&�pc�q�9";����J"$��_�J��;��y��&GC�lH���6���D<�ቭ��[�-�`r0��0��&��I��8Zly�!L��g=���sы9�9o�{Ym�QF�~A�E��5�
ɼZ��O�f�#W�gY��JcNߠ�S�@Lr(�t9��Q�����{��G�j�K]v����I�YBƪ`0����<u=7k��f�ar��E|���%Gܞ����0C�R̘�5~�.�J�A2�]G�Dn�:�_V��[L���`@���)�	5�M>P��B��ȞU��Rc���a���FO��%0�,���c��ӟp$��v��ף�U����|��H� ;S�9��`�B_}��%�u�Q�G+&Чg���6�8���Ħ�㷛�f !U2�@w��5~٭���Tp� xu_��s������H��m��N�?��O�ze)Pm`�$�[��5��{*�O��b��P��5���T����T�z3��\�L�°�j6=�K+@*N�ͼj�᷷Ng���g?k����N�v[,�a�+�xw��ߛ����g�Zj��Y4 8[��'�K�ꦊO?���(iE!�����H��ƁI�;���1�����3��6ᗘD��� $���sg��S�2S� �f��6\�8,����vJr
/U{��K�b����=��nE��ǣRL+��bVeLЌ�k�s)���s�>C��r�6���$�I�=��D�Ž��ե��u��q1�����
d�whp�����>�?Gy	S��x�8q2�NrLQ�P�I��!������
�~FӁ�Dt �BM��LW�,�X���弟�QA�q�l8>�l_IdZ����@m㽦*��)GFhD*3�7��N��(��u�����C] B��j������:�J�Oj�j�B~ ��Q=�i�wD�;tL*r�cA)�x= �-�w�ƫ�>ߐ�dJ��Z�)��w�[�lcd�ԁ9�.�W!,��3��4s�
�c����k7�T�%a�2,��WW�UbjB�l.�[����8�������H��0�Omt�n{>xU���g������I�6�o7�����2vH)&�"���T4�B��s��`�Z�(u��(; ��ϫ���LD5(�Wd�8�s�޺_6� �pg�aR

"����ƔV~(���[�}h|���cQԯK�v(��2�Ȏt� Ā����ѽ�H�Av�n0}(���zXgC���d��k0'G���!7J��hI�|����B��˒<��T)\@����
���[�#vy�Z�{��ܞ��(P�J�먆T2�ds-aP̑��"�iE�b%���3����!�.5w�A�?�R=|k�|�<mh���5�Җ��3��/���ƞJ�W"C�
N*���Y�1��Ua��/�|^{�x����,�����v�W�7���@<��+�<��m�Sp�����%՞�.�w�S�q�\rL3�}�t�i�9�����=��Ɵ�j�zRK��)�q��h>����1<������+n9򊓬��h��Zl��%�M�\�3����^"2�~�Xm�&b�@������;#��9�au�s��i���r����6>�����s:�Ґ�ԑ��4V|���%u�b�����?mO5Ӈ��v��X]dF�C�����z?Ԓ�6�!��!� %�t��U�}bj#M:�38G��U�P!��q�l�O�7�vkA+`�q:�����Մ�d�K;x^U�iP�j����!8��@��EΌ�g���`	�#�'�������>E�f��rݥ��{�\X������i�ް��[r�i�����c��\�v�S25X�֛ ��n�6�L�6M�.,8<!���!�C��,Z4|�O=�Aڞ�9�W7�9ٙP}�<3a-�U�?�nC��s1��/���D��=�����0��j�����\>��`B�$�.��� N!��h���3��a7�E���Zg	`<ٸ�����6|�J�\يK\b�*T��}����U�][�-�=��-�s8�M���4�
"�ss� �����٩�kĪ��E�t]�Ͳ��*D�w���%�?���d=?�4��9�zSpQ��uL�����T�<a6���JrX$��D3Z��D^�Y�fsIE�Ӎ�a���76GV��1�fi��!:/ _�0'���DS)F���B�y��?���ز�f!�Eƶ���8X�zW���C��ܟ�ˉe�ZHC��{U������B`�U;µM�Y�4�ZV�9SZXw��͠e��r�C:R���׻;9��=iDGn��#�X����Bqr��q$T�w���F;���Հ��� %���o8Y#���.]&�S@�-q>R�E]��{��.����B|��a�;��Z���� ��DBq����i�*g0�����I���2��J��}����xA�KR�� �4��:�)�l8����yU~!'M�f�ۈ#��z�ѻ�S����w��[�Ro�MGFH��R�G��9w́��:C�!L��W�.�h��f�ά@�c��@o|�����5�A0Ӫofa�Wz��/z�D}4b�T;ڣUr��"��10Yso�K:I�}�f�qX�Z��!�����TH��Zګ�B���c�4 ��	���Nm����FR:�~���_�����1��Y��Vn��7`}�l�^�I��M���eS=(��%@V�@2 L4���dv�p�̒�R#�"����L��aF�'�b�&���$�q��Ö(2Ih{,�I�'tĚx4����O�	���3ۊSpx����R�q_e�<�%C�#���,� :6�H��>���m�qy!�Sߊ���`�ozM�V�S��K1�"Mo<$7�@�-�΋h2�̺Kl�b#�oPC��� E��*��^���Μ���;���Ms*��X��,;�F� D�S�'q?�ѳLf������������sV����L�H?����t��]:Mәo_7��@~a��k�X�={)-1/��׏��QXӣ���7�LP�y *wq*��d�Fŭ��C��E���V�A[n�P7�m���]۠�}�i�Խ�ichk������[���=!�=���t��s;�Mvv������U��#�Go���+$T�6���P��᷾@@o<0oӭ���/E;��b��q!O�r[�km�|����o+zo�ַjmk� ������ �<+���O���y�
F���I�GMcb=�@O��L���3`n��v�J���[f���Y�*B�	;\kqC�&7�8���c3���cH>����ݔ~0?W�J�L~�j�}�7�4�y��"��0���:�A��;.��4Av+.�l/���(X���}i%ߘ�F�Q;үO�̤(�4x;9��A���2Ǌ���C��c⎏㾉d���+C�� \8��o>A��|��遯���a|�X��e�I1���Y���!�\�q�}��F���<h�lx���'��س �G+(ͫ�o�sHN�̸!�6z$?��jOi�x>�|������[#��Z��N�����H���������lDP�'�o��.�q��W�:���<d)^�C��CusD��4����s�&$��x�!���z ��uB˖��TU�)�	���x���N��jٚc!����a�6	+�BND�$�b�B��T6���Ċ�����jYvLI�q<�u���>�Z�z�t"f@�_;��0)�����q{�-����tt��y��C���l\��,���b�$�?qL���98Ia�@�g�&�DQ%���}���ѱij 冘�]p�vd��WR)�s���0n.�r�!������2�#9p4~�8,��ج����Zo("ӕ%��ʻ�5�a����)������[,���Th�h%-�.l����pK+�xޔ����GAN\mݫ;N�.���ì�3�1L������ZC�9���)z0�rZ|��U���I0��$1<J����+�w�t%-˗�=������Y���H����wp�20L�-��k����ި�a/h��&�4�[�#��l-%bx:	�̛�Wzl,S�66Wvחn|����H�{��N�!�	տ[�!��  �?w�&(�5u�_iH�y��Ww�Q+^��߷E�<�������E�d�!��z��B�Sy��)�I��I��)���|�;�!^�d�f��ߜl��m��>�l�,1�[�(m��N�=��Ţ��2�m�~&V�p�2������=�a��)SC9.y(����lLʄ��t ��H���5��t�zn|2�&NY���S�S�i��{R�Jk~�"�͡�}3�yD.~դ����K~���3y���]��9���+�qq��@�=@O�����-J�f)�������L�[L%[G��d9M� ����g��
��<Dؔp�+�t����o��`�ϸ>�+ �6۞Rs?�w�&�4z����Tiep���(3��� �V:�e�"=7I�f>S�c�R�\gI�|TC�{�;*�[��N�� @��,CqRA��z�Q�����GJ|;�>8�J������g2�xt����@&AJ��
��ԛ;�e�3����a�|������*z���?�ߖ����H��M)�M~l�)pԬo
".~����x�h�ضzv�;Lg7�@3��It��V6^v)n0m�����X�]	�"��Lϙ��? �/ˇ�3�3٨�mmڲ$L���%����d�6�l�^s',b7�G��ܑ���S��ƕI�2'a@ x�O�9e���*4�����Y;l�涫Kx<c'#D_�̓����te7���%�m�\�N-��|��T���<p���8�P�΍���J�7;�X�Ӹ��;Gl���C�ʕ^~YC+�7��������l�B��F#?ȭ��RB|�����gȳ&rI�D}�t]?��
�S�sdI��'��G��/XG�%�� �B�$�;Z�zи�|wO`M<�h�(��֭�Q9Y�]�Bw������=� �р�y��x�Sؒd�n1X���D�d]UZ��	9�6��J�b)���ip)��e��K��R���	s4�M^yc#��ϰ�9�iOڡ�k�CF��7�'��O`+�
B"#�̭�5�k������o"����p>��m�5�F�G�-�4P��!n���Kh9�=F��� FX� ��t��JX�\�^o �= �@�z��m����\�pwBxÀ9�1�9��������4jp�.���9+����l¶X�[V��E�0��pߞ�Ѱ�"��pw��ps��U�o:B
IoM��°�"���tx��6*����Ԟ�*�1Hu^�1���})(��,<��nl9�Ț�4�9�R`菭2Z�[���	ۈv7M��R�̰��C��]Z�[�q |z�-����d{vZ�"Ԟbϲ�<��V�R_��K�6Wm��Imd����S���OC��M[[����Q�1�ƄH�"%�@^
�6��*�t��!��|�� �@h��i�"y�r�ڕ�w�2>p5�o�bqY�"V��9oK��(?e4Kgr#�wM/3�Db�i���|~SAR�7��s���,L�g5FB��r��Q�T����H�)㿰�@a`o,$�Y0����yr-~S��4���"ֶ����W���N���3�����C⫱���"1H��t�-��jҬA�{�õΨ&@_�� y� 5���Gʁ�\+Mf�S_ц@��lg@�f����~\���,Gнs�Lt*0ka���đ��z�Tg�k�0=�uJ[v} Y�������5��@��7PR-\��긑�G�K��HU8��g�^l���U�Z���b��2�^G�{uV4f�"�T���]
��Uʽ~��'M�CY�w�C�3v���݄���B�(���I`�Q0�%�=�'^�[{�?0��F	^��f�+��/���k��n"��|ul��c=H~�\�m�aq��X�ȹ!��Ys�i�0�6ckv�?����Qz}z�(#:�u�n�8+<�����)ٵk����\w������q�'�rd�&~w�j�:���ȷ��1C3�lh!=�0��r���j�̒r^�1-<ffި%���@ǉ $�)ߕ�v�ã蓵v��5?|q��H@����j�%�28�X���<��6�5p�a��W���L�B�:3�8��^�(&��?AK���ёr�Ug��
hU�ϑ���&����`B�Ӣ��`k�Ϣ��=�V�3�����j@����`,�YC���ɼo���=�U.�WGR@��'bNX�e!��Ip�8��������o(����n]��l����n��4���2��Č�S&���q�|F9�a�����S�^I���l{�o�:]�sgP�W;2�;3�v�3�s2�N��9P�/��h8("T}�"��j��+�Ð�M�Q=�d,�Ǫ6�#��&����O�&�a�Vyx� ��JMZG?ʢɛ�	U�����Ņ�<�m��"�GME�q,	�}g�s%�0ql�a��uXf����.����,����Z���!�>�G� �$��)��W�tJs�R1���n���@`��[/
a�<e��_�Dڄ$�(G�j�lk�ˍ]� �g��'���=��
�cK������l��v@z�V'ܧ2����G�[���@p^��_���4�%e�����QW�%�&�}b-�U�s�@7�jT��c�y�ռ��S�hȀ:?O��;��[�ǜ*�^���{�I��7=9��ǆ�C=Iː��k3͉�Z�ݗD�֨ +����/1�e�&о]f��(��Kb���q�.k���yUS���
�KD��]eT�����Ѳ��vAK��P�`Ͱ��*��b&Ɵø9"Y7[���:|F�P�>]o�7$�ׅ�����?!�2HR
���N��Վ�܌fJ��!�U�h	�M,ă��=��o���0��㝥���sXL�6�E�D��r��j�$�e%� ��t!G�vN ����RQ�O!,ٞ�-~ݐ5��:ϋt�?�F�x�V�����ÉVc=w�+�����zO+�=�0>�&N�ĝ�}�7إ�85(����2��$N���[��}�/ʝ��=e�zƽ?(�p�9´�eH�D��r���?��x��n��SV�5�d�6�NĦi��~l��ic�q��^��aA����B�Hn$��J�ѣ�����x]1���`c��^�􅯜m��4! �̫Lw�M��w��N�rc��B���%MA�V��\0��iv�0`k�̘����|U�;�'�o/v*X�u��*~v����Is�nd���$��������g7��F�**�_ ���_"�E����o9��$	�`�>EY<P+񟩴���k���	@��zׄ>k�q	���H�;��o�"w�O���M�y�H���;��J���5�&��hr���gk�ߢ/4�Zw��`�e�-�I��eA�����uㅨp�c���D.an����.c�������S� �ПV�'����9�	�L���	��D&|�3
b�k��� J�cq�X{J��Zl+��>$�?�QOC�Aչq�lN�x��}^z�����T��j� �e�_ߔ
�f���2}L`M8�&▵��lF�~{J7("���K�5"�/��+2#�?�ً�C�#z����������:���M�t��	R�ڳ��7�Y,ysdY�i��[N'��bX�Q���/��+�!����[��O�4�G"���+������5�J%�'��TX�����XK�k|3�7F�H���1�E����=���;���� �݄�M��6�f���%�p�mn���k��S�I!&˔��
!�&�_z��r�=����͗	x�ZJ�0�s�,�.���Xq��3�j�Ͽ��p���Db�S�$�{AꙌ�/��6_�݀U|��-�3���T�����Q��\
-q�Ե���E\�y�cĉ�������sx�s����xo�4��$4Ǫ�bK� _�����f�j�4ƃ�<��1B�!��B�\��)�+VC��O��C$��i@(O��0c��d�B<�7WC�xKxӂ�w&��D��T蓈Q���&�&W����%-�ce�T�_���Ƅ3��Ah����	��^,&6bo�am!_�4���S��:� ��D���`��\���B�.���W���(�p�1~E>$�v����`�-���kb�6E��'>��w�^����ξIb��$ͧ(��z@oW 4�å���uLX�1p������ݱ�Sa��,�dϿ�9����Yʫ2Ă�7�}��9`��j�ð�>�Yэ���-YO	�JT�	;C�x�:݁�׊�y�W { ;��`]-�X�J�B�۳:Ɲ���s���n9�'G��ۢ��;���^Ǥ[E|�2�~��E���X���,��u8��z��<\l*�{�������P���4&�������1��a�����%\J�wF�K����t���{��ʨ�X��X��ϒ����j�&��~?��5��+���	�+Ю�%�f��(��_7���#|�9j�Ꮞq��D]M*|��� �l��J^qOs�f����%���ͧ�eG���ĴָK�}��bTd��C$����jǂVt�q5�ӁyN.)6�*y���cB��۰���X���t�[:t�D(\�Eu�z
Ѿ����Ӓ����n���$c�ň�e��R���+h#�f��@z��/�#�o�+�l���݄��eE�"b,����N'X�f�?p�tL�vF��@�C�C�~��� ��Q�:��Qe�[�ï�����r���.lQ�l谟y�*��&����.o�o����+�`���L�A�����jS��-�(N��|���|�xl6���	M]qB"X@U����H��ʟ�`��W��d����~�X�B�' ��[`��/l^��B��h��Y;���fooNK[�8��Cf��2t�����H7""5!D�{��x���@��>dW  N3yٙu]}��pÙ5&�B,���%H�*�����A�;�y����9��5߀��8�F+�iU�H�����$��J:u�����`�U�i�k��*��/���2R+GU��L���j2�B�YAk��@���`��V(jՉ��Tˍ��x�h��以7�ٙ���hVd,�8~{�da�
�������E��6gW`��ԡ�i5�}S�1Uh�+�緼�@�a��@{1橅��������$�^}�r�Ý�X(�x"�Ȫl!�ʵWP�]+��b�o��= B��M�G�2Kf��؞N��vՈ����wr��y���>�����.����Y�f�Q]���>
I�/��M��<���VRp�H��_E�g�p[Lq'�df��^v��p�0<Q��"�r����!s�.D��iܣ]Ѳ��2�w�4�h�p�eKϢ��hfn�+���i�ϖ���m���5L2�X��ƻΔ�� f�$8AH�e�E �8�P�:I|��̸�N[�M^U ������[e��-��vj1? �]����o���'`B�.UC'x2>V�s�_���7�c{�͘F�X�ƽ�"V�(�P$�}ܯ��Дx0'��|V(��P�1���<!��p�an7�I�#����R���U��Q~p&I�px!�#ԍ�_���h&<͉�Y!n-�tp��:�πJ]n9eL��e��8uN# ���e�c���z��q���]5k_q�,��{����c�p7�R#K��]��%<#/�Ƃ�ʔ�m��6z�څ�}�7�N���4�1u:��9u�N䦈A��2�^W!f4����x�c)F�d�ͼ��wb��;?X����\����ᬐ����I�`�S�Ă*�)/q�(��,um�d�� �+����9o��R���vG+�B<%#�^����	+���5ky?K��c9�W�l�L���&��z�0I�rUko8N�'?:���
��B@����B»m��4�F����x� bǤ�o���k��@��ژ�����ƳPH�6�5���܉
�����w� ���a�yqo\�h��!A��a�^܋M���OE�^����u��>����U�v7��O�dy8���oMhF��e.ϟi����N��EfX�	�H/��&���:6h	՜�yrRCe`݋gsj������bTiU��Sf�n�d��L��'h�GRf�ʹ�L��Vv��ȫ�7<��@]�a���)�4cD�sK���3'}Ҋ�2%r疿���^��Q�:U��=5@��%����U�������H�s�v���<���a�W��x��S/ܡBM4
4C�<�d�@Qa�͐�Ou���( ��=�w��&�7,D/��܎�e�+ҫb04�Ư�V�m������$�)l�GV-r���Uy�
��sѐd������OQ�m[���1����H*X�����~=�t��]�I)��c���-ztI��)��hot�[F���(ݖ�����<�x���o)I�g�15��o���)�]SW0��E�$ju�?�f���	H��5Kr�� L3g�Ud)<0�1VJ�M�u,���[U���t��;v��ܰB�7떮���,ќwv�.���;r��asU^�'4W����,���e��*1���U$��/Dˍ᪪�����V��W�Vc��"'\ib��0��̝�3 ���p.�c�zլ����{��=�B�z��崑��G��O��E,sAЙfX��S$�Ѷ���d|��hJ	��O7_�(0���z�	�i$�
��+�9��@x�ޞ���,'�ֻ�����xѕػ+����a�0�F�^4��_�q�ׇ���8O�Q�k�k_�7�����9[��,<Q�xg8��� �8K��pߥ��op�ߡ�f��n�@�Q�n�3[�����:���v��i��Ö#_ǂf�
H�KH1# �@�Ub���8�P!�`�`���\�K�U� `y�نF��m�q���5È�#I�V\}��W�����ȭŃ�~-�[#�w4u�A��4X�����1{n+c��	h�"(o����z�wn�?�x��Gݱ��{��/��#�G@&Ϸ�a� HG��Zp�@�m��G7r
?�=��J�'F����9O�\�C�ׅ�z����!��@w�GPW¸�a�pCf�	����J����:�j�P�l�=���t;<*)>	w��C�|)���\���P@��nZ�q�y3�&�X���������(d�H�ayP�g�!�ܠ�T0kt����kωA�����^M������y�$��m��>DK��xv�8X�5�\��������z���];�W�O!��m��G���7��|E��ҮI�R)������^R���w���h���
2���"��>��眺AF���P����r.�s�Ҋ�w�����wƄB�Z�.bIy�'�u��J���aHxy����o��4s�W2��v(F4�N��ph ��q �����iA��tkR3��#\]�FLI��:ȠP�	�d�}k��9����ug?5�9���_|<Bt���w�$7�I���0�E�:ۓ���*�ː]�-��V.Ү/B��\6�VX��o�K��,v�c9V�0����2�0�nj��%�����Y��؁�&.�����-�]MZ<���t��`�-�	9Ȃ3����Lz�ޞ����pMbl?u�O������[HW��f��=�_�Y���˧�!ϸ}���t#D�He�����4Y[��[�c�Sa�<pd�+��yh�N7q$n�h�ih5f��W���h@��G����[f/���'o��(�C����o���0J5e�M�&�>��Z�e�4��3�YDq)zq�p���w2_G��k�7G�������N	W��|ۏ��m�g#/^������ũK����cdQtAM��D���u�c�!G1.K�<�����<9ah��/1^�P_afÝ:��}��SD֤}Sǀ�4ʴ�`��c���:�ǶYC��v�c�2W�7���<���O�ܔ�W�þB��E��i����/]k��J׺�I���G �H3�֨��#|^R��N:�k�qmfw��}1���T0�;I��ZS����G�b�$�k�W�|���h�����cyQ�.R|E�z�`o�t�[��mg�GoE�CWJɠ��=�}�Z^���d���(4P8�dmZ%'�S2V*�9H癬J���z��N�	9�4�j�?!�<W�A�5���K@t	hCM>��*�Gz!�����4�����_ER�QlR���#bZ��ײޠ�K_�'k���9ބ� �_���p�t��� ��N���r �����c|ͻ�t��ʹQ6q%�0ݱ�{
��:IΕ�Sp�@��I�����gU��*tv���m:��A[��(j��IK��?o��7��j��n�I�A��a{�a͢cx<����Q�O��N��Ź7"�17ߴ����n�b�r�ґy��HL)�Ȣ�=��o^��2�`�;�F�7@�u)�)�r(vt��sJ<9�5s�3�RRB|����C_vZ፧55}9��$�'�3��M�e9;a�{�HKmo��L}��q�n�����07���W�s�)B�F��A�/�6s}�G�au�C����n]��=����,|���z��/ڒԴ΁J?�z�;H�D.�넞<�糪C�h�;�K�Ȥ��+��w�V��XEQ��f��Y�M]�4c���N�!�ƣ�2x��}��w��)ț�_��y�
{pS����v�B�4x�XXe�S
��vZ�5�����v�&����/a�G��H.�⺲��&�'�Z�b��bu��SV�*�bx�h��-�%��t����0��4)����.�����*�������D���P�V�5Ģ}����[yZ~,+�޾p �F2��ͧ���˯�rW�������<�I5�����;�d�#*�#�:[I�SM��1�m�բ�1.a�iߒ�H��푔���[J�g��9Ö�y������V�����~���#"����+�.��W��n�[�]R���'ʾo�^ٶ�Zu���j���J>fP�d-�}�*��vo?�ͽǏ�+��=f�=�ڇa��Ϩ}�<�#��^��>�yx��6�DQ����1+s�v1U�o�zW����*�9�ǃ��x�|�v�j�DO��a2b�.߫lE�w��7J��Q4�S�)o*+�x�D Z��rՖ����?`��M|j��n4Tm��C���<�OF��5pnh�ZPL!��w��QZ��
<�x0����ѾD���ʎ����j{ËnXL�-i�y�B��Q�Fp4a� ��7��E$��!\<���q��=�9}�j]��
�5:�\YJǧ�n��#�%�/]`�&2�P?l� ��R��Lo̧��>#�o� ������*1?&���}ϲ���>�;ߤ�5x|��35��BD4������Ûh\�ޜn0Px䍨��E��w��?������zp���Gk��~�(�D&m��o��ю�!w��	�l���[��>��2��O(�������ˈU�!�v@m�<�y�Z�KХT�Q���Z�Ӂ�b��8Ms(������)��Ù��R���ik��:^z��2ᙖq�
:*��;8�fQ��VFAT��7��v��THN�P�  �3����k����^н������-`J�[���E/���Vr���݂�jeW�����Bo�;0P�E�35\+�Sl��z�r��<�/e�ҝ���,�c���VS��;��/1��������g j7���mIh
��,���sKdB>,�&+�����98<67�^?�$�hg���iV���o�0dP���E=�5,n�� ~��l�g�?95��Y����|�� ��_�z�c��ŵ�q;��6���-�H�O�ю��珹���7n�&@�#
��FÒ���ptDH��p��_��k�n#e�Z�K��
�v8��Yr�0���]I��)G7�7���}	�|��v�0T���`�wbI��s�?N��2�Nj�ӥ��Bm˦SD���DqH}.��Mc����Y�U���T��
1��R�4I$��~�tyW��ݲ�&oWMH�+��Bd�Z%$�P^� ���hܖGMս�S��@*'�z���0��)T��ndK+���uL��5T�Y��՛HǶE#���)�g"��h�E��{h����p�iCn�Լ�{5 �h�Xj��uA�����.�I~��ĵ� ��ԭ�.�/�5]�1����[O����i,�˫#ֶj�����I)���܈-Т�9��2�$�A�����p�Y�W����<)>��T=s���T?Ṧآ�(�ɱW��Pp�w���t��z'+HEz�������1v���24^� (�G����H��;J����qx�M���4�6y��+.v5\<,P�aE/c�E	fh��2�0�H����SȯK�&c�>3��#T(�;]!�wd�����h���jaȒVm�fvyq\��$�϶�/�_���Ǐ��r�dk�I��{h����8>T�'�U>
t�><��tg`s��5���C3���ģ�i�a��%��)��ѧ�+9���븘����v�+�^WI
xŽ��\Ѹ���d�˺�+��^Ǳ�bO�0A�
�|�C�}p��&v-<�lv&��ǽ����+e&W�^�t����j���t,1�dЀ�;E��X��&ٖ|���os&b��p�a�<�$h�>����^��Pa�ć���"�z��H��cs���Q���oRݴ��ƛ��l���kϥP"�j�D���_J�>}�
Om�v	Dx�xd�ʚ
�7��6I�4]��ɒ*���Կ�%����~)%����xC���3�L9��Up��ݼ�,y��>�i<� ���wY&BAN�vmQ��h��4o��&�����D̗?�ݜ�e�7�7g��/ڹ��(��<�'�a�?��v��#��vTLZ���~��ؐ�*�Z�0\m��0�v�i���g@U�AZ���3Ѩف�$�����ԛwO�
�h'�� �x!.����b)��1s��h-|��(�ª�q�@�CأC��|RپZ]v�v��AsE���a!�vQW�⷗�d"�R�e�{�PQ��א���Ylp�Jސ�!�&�O��m�V`m4�R�R�'<�)���I�GC�[L�=�F���u5��`~1.٭�@��ܼU��*C�0�1s�)ɸ�YR9"�&����� ��E�ݘg�S޻K:n���	UgF��
�A�;��fp	gЬ�D�͑�֐��&�d���!sT���bbW������S�"��^����$��h#��d���k�>�F�tp�M"��s墟��5���5��x>��%��H�@���?U�eT�mF݄��=��Ta�:*5����wsMP㘆迁��3wk"]s0U�硯'��+���N�:�V%��u��č�hk��z��&�8�����`M��x��VC�|�W�8x�����M?�ݔ��oi���  ��c���W���B}|h���H��rH��y�V��w�j�ZЈ/(B�;#�b��-Vh�KU}RE/e5� _�*�썑!�=��ѵ�/xݝ�Ѕ�)fa�*WC��ا�M�̼����~��P��輰�:�D_|/��1���@KY%m��?[����'�)bn��U�s�b�YL�Y[g��j�S� -��sp��d~u+�j�� �%�����CZ�U�9��'3�U���o1P�|��kv`��	�&ث�9z�
5Hޔ˓fH�F�{�h�"3��O�|����U���h,n�׺���$��;�1�|�P�,�AG��3��HC�h�,�{z���ǍS%2��NZ����mi���+9(7MGi@l����в8�${�y.��#4��R}>nďcol��D; ^p~Ylm.#:d v��f�Q 5��}X�v��anq<s��Nv���%A�5���e��V�^��E%mkvh�FV�Ƙ�{��zi��a������O��y1X���	;�1�b����������N�.�V�-v��`0N`���c����� o�9:��YvF8K��Emg�0XH�K�
H��'�:%n���|j"_��Y���2VB��'��S_�<�5���=z�$�ȘȾb/4���~H�����_c*kGt�T�ƢR�2�7�_�m���VE�g��DDQ<7��Z��ةwҗe�/9���ѧBrC�yǶI��z(�-(W�S|,��ř"gP��p�J8-:|M�[r� ����������=���b�ݼ�1�P��u]�3C��qY/��#{���W����ϭ��w���PNމ���D?�
��q*��!u�:C�-�H���w�z�>f�8cҞD�m�(�0�h�	�z�7L��Φ��
�L����5��J{R����C���_�	3ʕz��D9�-;�5�ݛS��(ɋ[�x�^����}�>_�A�k��p�Z<X�L��Ao��'/�E��?Te�w�[�%��=��@Y,��O�4����ϞP�q�
F
��'o#5��ץ�G����v�Ar�_���hT ���b�E��������cJڼ����z1k��s�j���U�W�e�Y��)C����
9K"�5�˹��f���Q@4�l��Ȭ�5����KMn�;+J �*9,�z ���{�j���'�e�?tn
���Q2V��<m��l"�"Ǎ/K�B&o^ў���y�����A�_��mT�GhR�l�6}�5P��s����E� �u�.4:���@��r�����Zuc�*bS�B�k�H����c'Z�m4��M(n����6:ϛ��R]�aw��s2��ʘ)����ҡ!b)o�[Q�ۦ�	�g�� ��]F��X�Ɵ�Oy��j�6�V5�����V��-'� ���$��+�đ(�(�M(���$	���Y�AwUG���sm�����]jO�rkwb�CT�e�~9�׵Q�1*�n�U�@�C3>c͐gQ�^b��P}��C9����q��Kn�i�E�h�yWd�g�_�A��=iq���f DZp��v�l��q�Z�Y��q�r�,K�<��u�d�`:K����-D�IJ�e �Q���ʵ5��]⋲�?hF��a�]%6�n�aYh�p4��a����JR�g�ym�#+���$nZ�T�ج�	�7��HHh|�mk�m9�h����(�0C��(�8�Z�3J7Ǧ�4�y��EJ&�i�8�)0e�ON�-����
��jX]8�qO���k�TyNӌ�_^bC2��}xُ(q�z^*����\b(@�ha�@���"�ϣ%(k3ԃ6��Ϧ}�|���,Y? uK�p$�j��K�?�ıۅ�!�1��])��dFc��>ŤKsh{|S�'h�l{y P���:��
�\��s�Ϙ�C�NJc������N� A��v��c�`П�{��V�paI@wAw4��8WS��)rM�����*1N��y�܍\kMP�1���
4��y���߽j�t�3�w���>�d���lY n��������,?pr?�拪�&y �������4ݗ��?r�^�'�]�14X��ޅ!��@V9�P��)~�+�ru ӏ~Hʭ.�N]
Kk��Yp��U�mXR˙\mR����ԏ�~��@�CF���Z&�!<����p�ݍ��4~%&>%�O9��hi'��n��x�\(P�k�x��in�����i�1���gCA:�Vΰ����q��E�6�w�#�a�0?vC�Vf�����,�-1�9n᧻��l�^f���n�]Z���������!�~}"��$��"I��%�+ǝr9m&o�5�@q�d�s�����w"p�;���h�����6�+rܣ^��1;i��p}<����ꀷ�E��.j�\�iCC<����;�đ\��F���q�@��[�Pc/����=��G��Κ+	l ~q�&hL���ؗ� ��,�����k������0��j�`�k�AA�u�8�T������oQ�0���A���LtS��6gn螺Y�V� ���(�"�Px��5>�/��(Ύ<��K�nA58]"įo�If��0�ܵ!���Zk��O5���`��7v��:V[�	t��+����kp4����y�b�z����(��i�����p�H�#�|�`�׾��GXaE���)��{�	����S��f��=bVp�/[%����~i������<���$`�n�&R��#�z��@4&Y=o�b�#U�*�&q�򛌆V��}���`���vmC��7uSD6:�-������V�_����6Z�"���%��ft�s�*n�2��ݾT���)<�c�����`=&��>u�s	�P�%��M�ݍ"l�ĳS��q�4�$w�=�F���*r/�NKf��j�R6���a�Ɇ�J���o�L!�j?���D�kQy�0��)�ݙ)F[�v��( (���*/QQ����L�������鼖q♐(����z#����oq.��u��$�R���{g!�;�U~�^|84ͱ^`�!<�/:(�ɱN��/u���H���*؁z����p��4q�JW���<L�E^w!�@��ک�U����@B���hB�j@(��su������8j2$9ۧ����T^����0�*x\g|�uv�5��Z.�TmB�������;��,N�t؁^��y$0}��v���F�L�+��"3(�p�����ŞC�<7�9_��G=�ql����S��:�j�;�kU�c�"G$Θ|� �Uٰ�ۏ�C�[fk�rj`�Ǉ1hRD����Êz}d܎C��(E���+��`�-j+�!��K�}�$
���\BZ^uB�D�C1;��>��	P���5U��K\��#݂�b𴕆;F�Ab&N��r�`1�� t���YG�L��æEHq�v�gq�['��p�&g}^#����L:�,B�̒~N��s����W��C#����8J�����/O�~4_�\�e�h��i�L^,*�D�����q�Z���B��Dփ9��7���ץ~�X۵�d"��P)Y��]�x��!D�_�X���M���\���?�d6�XY�nq���V"#�7�'$6 �V��B��I(M2����e���l�p�Ҕ�;�5�C&���D2������]�vyQ<5Y���ðȪ��a�V����h_Ę+�>D �YR&Z5�x��*u�������xσ �mn[Zur���[���EP����@�T3l�J���6��rh��ڳO�4_�Hn*�A����y��&Ս�;v��R��VɊ����^� 7�_�ʙ2p+� �;(� iw�KU���n-$���q	O�Cq�,5A���fr��������#�\oa�"��˙�W�� �X�����(�d�[
���Xtr�R���6�b�����_��g�B��;̞�.?i��b�19�z\1����\��F�W��T�P���u�'VyF�k�.@�Z���D`nk�m�%�/~!}��J��[n_3���.�,s���?O��#�������(�u������La�
�/-�Ԍ��\��۠�t�S̦���qOͦ��/c+;n�}v_�d�V�)�nEP�9�@¥Y�z���o�%�/i -:	O�;B-�w�]SS���Wp��Ϯ�o���*a܉7��`���lcq
Dw}Cj�C q{��#��/��O.�-�f� D�m���Aw�;�wę�:nZ��Aփ�&9���ܘ�Xa咓z-��s� �"�.G�a�D᎟S��rH���_n���{�󯴵�]L�h���dn?�,8��X��Z��*��H��yv�	�\Iڌ)芗��v�͠b8QU�kx�m����pj��$��f�zS�<�;.#B��1�NeR*��"�����|G�<ҝ耊��q����LF$���Ё�a�h�M	���U+�r>�\��9�� �Zh��5��fI�����mJ$`�p�&ԪP�m��{5��g潑�_�4v���t-�z�4��MO�
�H�S��ƭCLl�>=�T盻�sp����&5&�W[-��Ѕ!6�q��d/e�Y�y;��g��� ��(�\k{꿇���ŏk����N%C�*�̓E�gʫȪ�"vuӠuP��7�]���&�T�>Y��~�� �Ԉ�|E�@�&j3@�҅�V��
�O���,�E e�l~%V�%�#���`�19�jd���u[ࠥn��6~l��}����l��G ��аW��oB@{�6�*��C���+��s���# ^��V�q�7	7*	5!h$��J;���Z��7Mwُ�Ob���A7C�{ayu?��Y�;u�R�l\��V�+Z�&���%"l#il���܉I�Ķ+�H�.��v�׹C���Đ�N����֔�
���g4��Q�q��J]��A=u�[J��3PKw�E*��1ə���y�>X�ح�TO�A1��� S]��i�H�'McI�r7��0�O�-c�MT������=�.F%x�F��6�C�yQ+϶&޳�4GZ�O���tҠFDCj�$E�ۂ�:���!�Ҭ�I��X*�%��4�7%N(,�ۑ7�D�B��y��ȡ���O�V��vӛ���x?�l�#�}�����,��L�퓃�]~G�<?��	���Ҫ��]`�M�UAD��va�}8?��D��t(�3W�^��$W�
B֬~�3L��Y~��*���vz�!����,v+$`�]�qJnOs��!i���|��Y�ߩ��Y����y����JNe
.lY�U��#�a��
E��GFg-c��\֪���Lޏ���p\jL	b�v���E�oyz����c�Წ$b��9�e���AQǌ��@q�8�o;%��Fݼ�����8b���[���;�=�/�u�>v�]��-��c}+�ݪn�v�e�R�U0X�ϊM+_0���P���Oxt�Y��]�����k?�6�h�NԈsh��o����5pD��b��� b�4��8*ȟ�.����=q��u��p��h����M��q���O9"E&���Zg�F�~ǿ�3_n7=J�ċ������^��j����ڦ�=;q'9�&~[��fFE��<�xh,�z���fDGV��Z&�Ùʢ�,�cg˧��ov|B��3��%AA@S>B1��� �7@�61atT"�M�|�y�斸a�Ƣ�*,D)����m&V�O���<%��� o�����Š���$;	�š��~��TtuUa���h��?���dr�LŬD^���iA�D�.s'̮1§z鐩5��~t�E���q#M�ARl�ɹ�X*�`��K�Nh���1������S�C�Mk:��H�V|�
��k,��:��޸��n�n)�s�v�r�o� 	A�6���q1%��d�j
��:�I_��_-n�g\��#'r����i�������ڴ�ҊQ_0^M��[��݅x��'�GS� |>����J�,8���!�����p���F�5	���@��9i6��2��<�%X�eHF�,��^ݸ���
Rw����(�e���B����v�������jQ��Hl,�zp߽�Ğ{3*�h�w���V)L���n��E����w~� iWZ8Ц�C�uY�.r�Q#4X����{w�M�!��J ̞t�����%�KTck�^hc�0�3?�J��2 ��U�&�����t�Nb�rQxҁ�wQ�9M ���*�A�n6nL�o>t[�,�Z!�e&�����ǽ�@]U�O�j�`!��q�Hs (pN�w�&�Հ1*`���N%�$����]�����Ml���҉�j��&���"B��J`1u�o�����\�#��a�ɘ�@2������Kqa��,�3*�ͳ_ �Xp�	*��$��z2�1���?���Ȇ�>��B�c�=��m��gB��Q��,��0����?&�>�����(�����;K�s�v~}�{�q�D?g5��J"�� �V��R����-�|�,��+��7W�JA�������s
:O@n�/<��<�����J�G�˝� ��F6[m=�]�B�&Q��c1`��SW���6w4�OH򹘊2���Mk��Q�B�F�0jk`t`*VF�z/�W6q����g)�W�0&g�,_��b�_�~�N{u��a�@P*M�b�~��F��8M'�_6<�b<`�ּ��a)�ir�(ʀԢl����~�Vq������������9���o�B�bq���I�5ze��:��k���T���}��kΧ�����p񯠳[Z.�М\�3_Ep&�T]�uҠ߾�)z���L�4!*�O�]���N%�e�5]�䭫i���!m93y��4�S�U��ς���"Y'�|�x+�ϡ�g�����}��WG�_��w�UjWuO(ck�ݞ9:��7�H�6\hn���������m�s��𰄀dG�܃��k�2��2�zk:���K�����Tz]k����1�>k�*9Ê�}��[L�Ϥ�KA���
ƀ�a㢦��=�s3Wxo��,����i�U˙F�ܓ��.�6,1�$_=�=��`�-�cy���T;��G��*�֮"�	�,W蟂A|���P�_�A�+D���+�����U'�Zc����tuoQ�2����:�.dmYp�/@������ܧvpd!��Щ�v5��w���iK���0}��9�!�+z�Q�����DzxX3M�L�6;upRG�#F�(�|��z���Ȏ��Xw�Whh�8@���+6�$>�j����0�i<�n��j��n���ڒ�*�ݝB����aٱ��P�jr�����(T�[�f�%^+c�xC�׈���ee!&�P��o�&�y,ƞ��d�{A����ן�l�<��3לP�������_<��܉���	��}=�*��ȵ����x��oM�WZ�L��zpH�.�d�����ww5Ck����ʪR�c]�IJ����4�D��ܷ*!M>B�$�-,Uz�y����Ǧ��?9�}gU�Ϡ�(ti0�q�����F圕գ�Ύ|�N����|w���8�F�s���Lkb?����Hg������y���iN����i4��L�"�5[���sފ?s	}� �Fe*�
Z��k���Q���$0��٠�\v�\ s��}���t��HeQy�^��Ԝ�1ƅ����#�U4� ?�PYL�y��l���܍�L�+b����N����"�C;�c$Q���Y����%,&띒�y)#��$��I�
)�y]��&�!,��!�0j���"H�ߏ(D��{\~�s�6k�֟�bU�j~;���Xm5b�-�M�~B����>`Jo���1�6@��Ss�F�/�q��0�z�D��^�:�����	1�F���m�s
��ҟ!�A�O�fSư`���Wf@!;k4��u'˘�_� �,�x�/5B4��6����� #D�	��N�[uSP�	;�g�b�ݲj�)^�?bN�s�^�����H.�����C�]����F˖�懶�����f����H4HE������V�1ۇ�e����֢�o	T>Zm�;�=��^;��>'F\>�]���|@����m]��-�8�����;�j������/f�9n�q�OH�����<"#��`��kx��6B�0=_��u&P��ʢ��_��������D���|�E"���^����
��
kC!���B��?a�8�k��N�ǹ��yw ���ʢ�e�n&��Ⱥ�����{�ٺ����Ѕ!�$Y��3�^;����:.�
x�m�o��$˳U���o	_���^�rjk]�!���t�n���i��`���<���ʉEİ�M������ώ2��@��K�c�2Y�Н�B�]�4�Fk���!Ś�P�x0=����7�D��-=! ���џ}�LI��vA:����p�x�5�f�w)��t������U������rg/	�j.�e�Ý��jP�A�U�)#��k?��#�Œ!)X�%l�ߊ�\zVⶑ�DS��d�����9���L:��_];g����җ`����3���`XDw�)�졈�rE�p��GѻO�d]���F;;��Ђ���,��J�ϥ����X<~�]���F����d�͛e	f�a�5�(W���y���b�MƑ��٠�UZ!|z�� 8h�cc��.1?��-}����4�`@�D,��eb�X��Z��X����Զ����$�}q��C$�Mt�#->*�x�Y����틻��?���:O1�Fa�}��2�հ˝���X�¸�:0�|��}��/���l�8ڇ��(�iK|�-w�Ż"?N�β�%�ۭ�WGQ-��+��y���b$�F�P�4q��)Ѣ6g��߃�7�a���ҏ�>u����̸U�tBv��#?����)�#?ɂ�iwv�N��������*��^+����Gf���]��)`�G#�gM�|��m������� �E�oƺG�u�bN#S��>�>�G�1�>Pn��o��]������儛v�VRTY��p9�k7x��sA+=�Zg�o��<������ӓv���C��	|[|��
�	����Ȟ~�~�M��y�,���#փn�6��d�8����P�"�&�J�УBԍOm�7��tՅC����&D�9l���!I���%�������tp��Oc5��ke�p��!��|\��I��4֟S� �V�"� ����-�P�H~�{��"�2�_��4kf��ӈb��U����s��K&O,x�,�
Qu-c�&"m�1C����-ވ6�8�rA�
7�'�|�T	��ށ�;5h�K�n.eU:p��=J��+��1�"����k���s��|�T$<сd')���M�2���C�B <�Ռ�P������5�}f~-zW�U��v7"�|i����wJ�Ai�p�E��}D�;
#?�h�^��"H"� �N�B��6<J��ܩ��#�daIy���'�7Cϡ��|�`@&<��\��������(��.���y�@[^QWW�T�J��|(��;��-?��B0�BQ*3Y�ҽa?{�:YOqXG���f|�k�f�UǤL�,�8��$�C�y�+d̟R�~'�II�Q�R�p�Mü�١��KП�FFT�+���j�|ےd�p�����jⵔ�v���hp���n�$'

G.�Ϛ���7A��x�&XӞ�Y��J�B���+>��Ε ]�V�%��r�?k�Cq��8�Q~�dΠQ�f���=��N��ql�ui�89qi�\- �)��	��wؿ1 å%'=��1k���_���*�E9�V���>3��,�YM�D��B����:5���)�b:i��(u��t��s7�����fj�X��,�����ؐ���wJ���c]#qxׄ ��4���-�~M��Քc�9��5��{�6	��"�7��PK�̿�r��W�*�tf��/$�:��N4 4�g���'�}/ N�S��3�����3yq�鸟͆t���94�����*of�q��bM�<>�ap9˜����+��(WO~tA����D�A�z��y�Ze�2�Z,-�����_1MҒ-��NpZآ��I��	��h���&�E_1ŷ�	/������#DRHd4��\�	c[�ql9����O������E�j^��+�&6��I,�n�Y�bX����rۯ�	��aB~ Ir܆W����۴��\���M�DT�Q�,�n��
�їnt�9�v�6�����ו���b��w�iN���޺��l��)�R�CűK����`�g���f7u�O�o��޹}</vxz�T�>h�c��#wc�!�mTi���c�����@�Nwi�HA-���|C ���t�ǌ���y�v�~*(�U��X
�h1?UӼBw�Y�k�����:Y�7a����L����"�0L�,��QQi�ėe�2�Py��o��
ZѱEŗ����{�#60m}C��bQ]�=�\]So�Bk��������Z��Jzޯ��cІ	Y����b^b�~�XQ�'Rh������V�#��y�z\30?���w$8D�ʓ!T �N�g>M#y=�{Z̒,�)يG.��������֟x��1@xe;'��*:���Μ�ŝ!��4�
��QN'��iCHч
&P3���%� �/�f��}�df�%� nb��m����~�П�1�6��j�?u�;��l�<:D&�6)-����=_��q���<L�s8:��(+�����gpo�T�����q� �e`4�(�a�d��f��.�Bp�j/�燌*�����A<."Z,bGmo�@r;{AR$�"�N���)PƴBtZs��Ċw���|�+�t�k��"F� '��7Y�E+���p��fS���I�4c� ��,V#����h��gZ�y>��[�$�~j��|�&�u[�S3�$�|3S�Š�yG���ho��o[n6:���7f��3,K�5�X�	]_�,�E�+�,M���P4�I�<N�iQ,3�E*kLel;�՞jU����9 ��z�6�`*S�]aﴕIqu*�c�3s�ל�_<�Ap}c��`�E@��`X�2��+p�������K�XJ�4v�ب���kfA�Ѧ=���m�]�`J�%�c�V���l�������d�Mr�a�f>B��FsIvz���[��� ��� ����"<K�]�(x�|"�>� R������1͂���������`7{���c��N}��Z�`���	PsP:�qEPh������.��{+���M�zY�Gjx�-[.�V�s���`yCkJְ��̾���X� <2@*NAe4|.p)u�9��}^��2���F����y�9�qP{K��#7q� Z�#����0?�GzZ@N��	W��Hc������qD�'�*+���f-#�	�;�N�0+VDK�u%���=a�`���M�*��5�xޗx�e7�{WE���Z�c����ܚ0L�U~q���#9�Xz�-�'�3	��Ժ�m�hĕF쟬��Uds��1�]�#l-�a�X>� ��A�6<���]U�d��bGR/#e�{�R3���A#� �#(�[.h���^obL�MS�c����)c��a9�T�&_F�b���$f�ӂ���cH��z��_O�
�	�e�tOmZ.Z8v8�ˤ��	w]���)c���|����U%����LAX�	����*�u�:7��]�8|�ZL+���䭺!�b��JȌ��H�@��BIǖ�� &d�����ZD tyT��g��*jQ�Ȧ���f庅��!h�t�sI�$��0&Y�9��D�v@��BY1m�, zie�;��\�?��򀍕k�{UO&l��ʌ��$�6�x��?�JgK. ���փ	s�H�;	�3lQ����Oݮڛ}��,�m�j"-�S��.����׷hJ��&4@�A��Ͼ'��=?�i�ߩ��	���S��wCS��j}D�w��=�0�֔��F�:��W�V�&�����WS��H���tz�5�w�'������F��8ņ�~�C"��Gԝ�/";*� g�ƵF(����%�A�گr��B�J����7�l��z�=ga��Q��h	�N%�V�n�i4X�����H�Zn�v_�~�!�bZ�r5/��'�Zě��`.�E�@	O�Q�n��I�~.g�D�,������@�2Z	�j��e�}b�88e���cD�V�b�=��Zz�g���k��C��[�	�S��,���E�m�,��N����������$�7��|P�Rld7����fm5D�l����x*�{OT;���vq���4��{�3���Z�����I_�mSt��>Jx�%
a�3��-EN_T�fȼ��w�9���|�g�T:z,4x�=�Ŋ|��vp
l�5MV��jefW��A��Dx�NI��\�f${M���_��
����[+Ny��9��{�������M(Ǧ>jY	�l�*��* pO�.ʋ���Fo����-�1�P��`��<!r�N�·H̦����7�m#͹=��D
��Ӻ����d��F�;�ʞGW:(Q��m�,��>ߑ�ޱ�`[�m��}
~<`>[y�G��,B�P�{ҹ�F�W�S��-�X?�.��0��a��C��0�D���$������zVq&B�B�f����910oq�hf����;Zɂ¬פ��L"b�Y ٴq!�m�ԭť9��F���;b���J����Se�ת���&=����[kS�b4�%J+�� B@!����	�.9Gk��Q���sm�X"09f�u~���]�(8����p�M��Ń�ƍ�� �Y����:b	���%ƹ5�)9���Ppg/r��=�mq�A��ܬ$Q!9� �^���ªl6�S�8��02����@��>i�^��ܱFWf-��6j��-���U�����3��yE#g��2���n�@���-���S�p���è��b����>�Y���'��R��f�V!�D�ͼ���=�>r�����KI����8�ѵ��!��R�<�g_\'��܎�E3ݘ��d�*b\}���e�@ea�`����17|� UF�P���xg�����1�ul��]�I�İF�$��{w ~v^b?��V�=E�!�ն\��Q��ߺ�=��:{���H&�0� � ��t�������R�4�Tȳ��_�hS}��i���}I|dA���ʶ����%���.-�x sg���N�����:./߯�L�@�	6?�4oټwF��Q��ӡ��ʕr�f\��S&V`K,!���},/t���r<⤈l���=�9~`�2��O�"��o�	��PM�Jb�r��&�UgTT`�h-}�e#�֙�I�:)�sU(n\����3���,Z�ʼ��iO6�y���C�lm���V��/�^�X�g�* �(Ee�N7rk���{�aXzUS��Z��b����1�	M�B\W�G�LO�/�P^��2&L+8.�'Oʷn�XvR1<��z���B�R����AĨ�,�
:�r�I<���z��/�:q§C���ȑe�ľ� �F��Oʝ�]�$9�}ل!�4C��p�RM]�2�T�!Z�8<��׶d����Gb�������S+�V��l�G�Q}�q1dTw|x�n�Q��Q�B��-�,����^� |
�9De�+H��^�(�����1'�nX��c@TЊگ!Ό;Һ�?�1pE�m�Od2+e¬"�ڹ�/���'�=JaW�� T鼑UN��p��{�b$g �~�@6��{&膱�=�N���Fd�'�D�6DA�J�)/�{�܁k�\3�'�jta��_��O�-a<c	��Q`��D�Vfظ=��������o�n�D�#�5ݥ��6Y8�,z�Q)?���K�N��b����lG�|���9a�i:*n`��1�,��'!�(�g�����}s~Ʊ4yEJt�0c*�����I��uĩ3>!g٭��X���G���}ڮ�O��u��?c�;%�"��M����h��/�B��o� ˩>K���t$͂r�30H�(5�wH'Y3��h�,����ێ[n�t���D?5��C܃#�W�J}�zD�az��[�#;<J����/�����6�R�ta�?�dnt�L�Pi��F��ڑx�g�w��'�2��&��U�n�fa��M2��TN�?"d�M�	�)���K�Àb�;�Ӣ��KYDT����E���$�T�袪sզ�u��ӄ��*"��P���-c����^�~o��2��gA�lT��)�G�RA�HVX��Q��"�&,Ky#��B1e�d����YIY���>��^�X!=�q�.�K�'0�����g�]���醯��f��Y�CFL��1�P�~v,��V]Y�]�w��ҏ�́�s��m�U�9SD����f������L��3����m\$�(��B�hjs��1��p˳���bD�]��T�9[/h�l�;��sy�C��}{QND�	�[H_���}�CG��J\јqxa�� /j'��5}�#��W	�e���h��`F���7��z2��4 �*�F�"s�.�Q��2�Kg��^P}PKSk5�KR묥]%��xm�xlv�vB�%<�<�ȇ���V	���0[��iƅ��.d
��&����M���-�^o}����Iӱ*�?f��b�m3�����,8}��c$v�IX��U��k�`���i�q]JMz[��C?�i����។�^�,p*�b0#��g�-!3���N��)՘���V^�n&��N!��?�=	�!��&6�9����$��J��Km �A�p
;���DB���K/�V|"�ne�X���̦Yj�B�=�j�t�[.W��&�ҩ���}v2L�.���J��W,I(l�mﶂl��[k�}�͈e��;H8�;��x�w��CA�4Z��N^���op�?�b������0��~C��t��U��:��P��#>����b�53���e� >/n-+Q��Y���{&E�`8��5�O���5�pr7��J�O�p�J�\��ݾ��-��Ph(�ت�O� ���47$s��*��Ў�uE��8 �΋+�-�">T���A.��l�F(&H�в��>��l���'5����#"��er�853�� ��(zȞ�����y	�N�c���ό$��'/���;�w]�08����$/������d��p|��[�c@�`��~	;���������iaS|���R��`"���~gô܈��j����AjR\�	�d�
W�F�#L�Ϧ.+[%�����:���חA����@s8�:�����������	mZ�c���J���Z���d\u-G��{֠�0x�x7B2��W�J�"�\E�As�c�Ϋ��"3n�ե`���Pcr��p�C��W��x�V,瞀$���0$���{�tA,U���37]�ыDd̎����wM�.k��Hw7�M�/N���bԫߣT�*Ԏ&��ڤi���}\�+�Ъ���#GЗD�'����t�n�����ȫ

��.�#=�1,��h,NֵV�ԗ9��'�H`:<�;��I�~6!�Pu������{�{6 ��p�_��JW`�8��M�+��_�_���'XgkX�?��x��&��աG��^��h����.e :�]3L�\��+��4�_��7�	��T�es��
bb���"嚡  �x�6A�C=�'�FP�
Q�
�F!{R��p9�EH�K�\u,7�39y_���Mƒ�R�A ݯ8P�>_���D�h6��9�
<���< ��tXs
��@${�)9��Е6����/VLtq	�:��Y`��| +wឫ[��x�'zM͑#�(u�9��}���@h����Icx���]|�rn�=��-Πㅹ���(�y]�R����س�c�c��՝Y�wO��4��#���̏���G�*�ƅ&��U��Y*�E6���_-�������'Se^�t�x(��  4��(�:��̴��`�����GU�#:��_�©BZ���b��4��@C�XZNg�ThPLׯ��2���GT?�9g#�&THd�<ڼZ������l�`�->��J�r�o�ƜCX�����zm:��\��]��1�#5Ke��3R���Ѩ�ˀ�����E������~p�1t�-}�l�9�z�A3{u��/X��"���ٰ��pha��{[u>J��3T��|�3�V�1�18�ӎ�|1���Jt�>F�Z�Ó���S������xHd�ޫ���;���5�T�S'Z�dk��� u)˺v���s(�.��K��+r�0n��1z{����'0H<�.Z�/vi8bp���7-��Ĉ�}ͥ�{<PYN�N�T���Q��4|j	E#�����HY���B��9 �Q��H�/!1�S�{{O��1瓙Mu���dL������6;6G�A�ᫎ R�W" �R�A��\����1��S�&2�gs�h(=�$�x��M�za�����'S�bM�p>-��Q&�#vA�ܽ\��{蠢��x��V�6�r��B��c�SB�	ӍOG�X�g��<C/.)��R���/'�aU1�a�
z�f4��Y����T P�,���3P�k�s�YCHk���x$)ُ���ҝ�^��B~=�?��:N�G������<P��n�g{�	�B;ү�7��>����O�5dS�R$��T��ή�'n���v#�Yּ�\�N�b_(�Վy6w#���3a�y��;���O�
�@��FA���U ��Q��P2�U^q��e��`m/�,�9WK�Q�!��2s�>LؤX{��Q0��_�B���y,�8�:�#�J�=���\���_ȫ鈫��m��R���H�+�u�����7��#�����|Q��+S�Hu��B���YxN����v���*���?������@W[P�%�83�{ݫ	��Ќ��N�\�È�QXt�h.Z�=�x���\�v٠���._E�h/�@&�=N���K�W�d8B�p��@+�!`LL:-���H�^@�F"T��E��`���ޞs��SO�91NԬ��_w����rq���.�q]=��\���ux�����F��jFwHl��-.	.���[�8�?)�q��L�eIMrw��?��y���"-����U�	�Ģ�����@o���(H�am#��,���[ƐL�l'q%h�(�w539�\<o�F T����O�m���{.M2�Q)���-W�����O��5袣�O�b�y�$�>M7 �>���Sip����n˼���ң�Q��1^�7!ܮ�v�G�IˤR���U2�L����ԃ��їU�o�r�t)��v�R���6$'�����1j�U/ ��X�._��L��C��ь�5��~��?MtvI7�~��^�U��+>wILW���	*�:O���z7�������08�]"����f�7��*;�?2MS�x����@W��r5�d�����)�������n���e�=�Ȯ-rw*��S,=_<�6�0�tn�����L�(vT}��z	���Zpn�R9�<P���%?�0���0 ��TM��ս%�2�>n߄���&I��jx�� ,��*.��P0��N�=Ix`M\�?)2�r|( ��eO�_u�O�y��=�£�ТJ���ޯA<,R�&�^��v�nu}K_H�mr�09�I?m�L��/�kMOˀ2�ڪe4]�s�lJ���PX* 5e�j+܁������ea���߬^0E(��8d�pm
���iIQ.N�[�ʎ)�M�BLɔ���������ULIJ_�����>1���Gr�}7�Gc���85����/E��)%�X�چ$e�Ř�ee>�Z�����$�=BƄ�}���K
�����)�]MVD�e
�M;ǖQL˖�w�ψ��S=Sx烡�E4f O�� cت/�+�/5z��A�>���TU�ѿ�S{-�{�J��P {����"��]V�9&e����2Ν�%�p o�S�n8
��WLy�����\��|�s�~[�KyӒ"�Rl8�s���9�=����C�sZ���r=�_�k��š�i���Y���Z�ytHf�y�E�kŃ�ȒA@^]�H"
 ڜ/X�Y|6��\�`1�&��k^���T��wԚu�-�g�t�GlN�j��������O�ݿ0#����~�fQj�.e����O�'�٪�B$���HݙFY� 
��>���Ȱ��H��O'��S
�)0�q	�D�6{s~�TRzɓ�M��� ^�����^&��V��#�v��[��ي��P~��>|��9ʓ#
FS����}�GG��8������.õ�\�j���5˂�4ܴ�X���3{��n�g����)�h�	T�9�6������l�^���\�5�f�s5�\�M�b�Q]�S���^[QB�l@w2F\ѹh&ԳےB*�Z��#]s����x�����5�B)��Y���]M�CY^&&��6��N���42�Ɠ㋰tW��#�)g�}ށh���E[*�EF��֬��\v���toiԟ/��T�m�&����ȡ���s�}���������B������K)'i�zW��T��`z��'��N�7�77�r�.������v�O��� l��/x��]�M��&I��`�z!{�۟5/�`�)���mg�s0|�uf���u9�#�8�g��:��Mi}Ҽ�e�-'��N�����|w�_fD�s"�a>�^z)�F�pPf|�3W!��NӤ���sb1�R�ʧ��ɢ(b�y.~�a�����wu�	�A\}��D��H�%D������[ȯ}�J���8}��K�пe[�����Ǟ+���xQS�����J�P�hf��^*T3�w�X9�,<�r!y�{I�]�����aN���	=Gck��X��~T~��B��6*l�����JZu[�ZF۸��2��Հm�9g��j��Rr{�Ww���&L�݊���!�Vz�iw���[���`�j�x��M(�7KG,p�r��IQ�:*o\M����ͭo�A�z��j<�?~���j�j˂� ,����]��7DO5r͋�vB��Y�����-=C�Q����Dy_0Q)̤`'�3!"YC�4�)��Q��1��� �@�Z�$��eK��Dq"KI�/��L���D<�E֍�"��U��4�ZO����ohhҋˬ�u�E�8F����G��7����2��T?hLT�x�}M���J��_l�R�\;����{��6n�_'�/|I��L�㿌<��l:m���6��'�b^��%5�L�o.��"d�?�����&Bӟ�����<��|�~�ͧ4�ҝӸ�'ޚ\��Ӱf�*8�>�o��Ԋ�Y9@�7Rb+B{�u�ݶi�l�WU�o�V�����%������G���{b$&Zݾ���q���h���ҵo������T;��q&1��������KJ:�
�!(\Br�7_�1h�[u
�Y�j݆�t�����vC�W�#�f`�
=��Y��ɐK]�q��Z?���TdO�M���͵5~%�Z�O�8U��K��l������d��LtD����G�^Z�<��T+�`�Ѕ�e(e�O�5��\\�'�h)b�_�^�|��c���`y��#D�;
4)�W\[��kR_g��U��'Pj�W�6C ������Ol��X�R���S�#&���_z�~fهAcͬ(��ڰ�g'v0A�	�D��KH�GO��g�P�0���&W�;�v(�l]ʶ���Gg?��ۆ�{W�f�
�ƠL/���4���f�>�J���V�;(����B�(nuFE	��q���Y�݀mZ\���oF��ӕ�i�mx^ޑ���	�M��_gt �=�(���L��gx��k�v��}Qt~��x�C�H\Gئ��@�S�A����(��d��I�\�zdI���u4QW<}1#���H����Mu.:)D��-�&N_�A��lQQ���C�D?~�&@e�Y��}�_I���o�}�.���������1��0��@'�!�ldx�(S.�6hlcJ�y�DG�b��{����`j�K��Ŵ��²[��� ��e���B��"4�w~ҭ<�cl�<�����=V��x�� <�>ϑ�L�/����]����zz�y��Պ�4�#U�i#2�ӻ�ˇV�O��\�`*�Nx�[̀��jl�a���E��'\���xh�3���c���f��Iڻ�
Q/
:��1P��/��f��q z�� בǁέ�=��\��+���Y�1��7zd���=��zR�d��u������ìOFcr�����6+ ��a�OL������
�Z�]d���@����f�/�fܒ�����F�`��� O�2s�vp���A��x��w�(1���=D����p�O��a�����UWVm����'��t;�5��fx
��}���*toKRj01�/&���S���%^��ROX��S��m�m�~/U�>����e&w�>+�2��u��uU��B��0��7л35��Z�ȳDR�:�s������~� 6uJ�l�l`��̱6��{w�e*�N��qР@�r�1H�����h�9�;dSt�����1�`؉���Á0��� �6�B9��9�p�쭩w�#��lԷ�50j���m�;��ჿ<PW��_��ߝȪ�F7�}c,��j������X��������I�˅6�e��)�n�A�P�?�EF�X��Q���t5Ƙ�S���ȇ�2�Q1J��ͪ@{��@�q�~<2��mZ��&\.�>ۙ����Q8�і��G�~ap��$%z	��KA .� ��Z�egfP +m5���i���!��sklZS�M#�m�YvKH8��H�©j�u����-�ַ���������6�N���*qǔ&�me85̓���M��.Gm���;�9s�~�P�$K���O��p3���sͷ�碈���[Z��V)q��\��������&���z?����9�b!L�cw�!��}bP���j�hx*����x-F���v|B�m���4�U�N�wဤ<O'�'�oa�"��|4I�WvMP>j�)�Z����	qjŴ����'�fA�1r5ړ�uɦ�[����Ғܕv��i��h���^��1(�={!p�k#�.Aw�V/ݐv\��s�A�׮&}�4�oRgｫ��i�G��E�b����Ƿ��/��>qr�kwu7H�0K�_�2�ZFLi��m�[F���[��8	�� �O����N �V��'1��s��%�.�5�#�Cǆ�M���F�
�t���"-'\� �Qj�
�%h��FX��b��j|�\WZ]~�/��*V�$��˾�f�]��
pptG�̪
>�����26�O�n�J�M�����6Ax�i�%�~A5N4g�s�p�鷜�e���lÀt��ף�C=����6����~��u���ݔ~>ʓS�%��ԌS��\�Z���Ƞ���*@���J#��,�?{aSf�~f�i�.�����1l��Dg��E�j��;ptk'�l�/��Xp��diO��q���d�.�aFC=��TM�!7�X�y��Z�_���#�{j�]wO����'R�	��0//��4�W�ĭd���V�F 5G��k��e��]l����{ �^l�I�����&1>�ٕd8�S���^@�Ip͞�Tn����Gbܯ��c�B=��2;���v��S����KA�`�e���ʣ&
�x���X���ᾊ��+l Thj�s�{���,�Uo����'v�Т�� ���b�=Jo��a�_���RTp��	�cLO�;f̀�f���`�P��� �(����_�lݹYU�Z05�yz� �g$xe�~�ofm����Su@ٵyq�ǟ��9�s/��!Q'�ɡ�C��F xhz�@츄��B�Q"��![/�����E!�8�C{�#�*58�R��Cm`s��k�j����t�I_�d�C?�vĕ��"�jL���w�D5��
Kp��@�X�=��nO6_E��&ϰ	��cs)SB�F]9��*���v����f�j��:�OV-Ap��Jk|��1�'+�������u�xG�10�����?M^kF;z�j�.!�
e��������C#e�a�7!��ss������:oq�y&F�h���͠�Af���!n|LY���A}h�
�#�UF�"�v)�s�cNp&�.��}�/0��c��Q�zP�m%_������'q;
i/{��X��_�<xP�e�Z�) eڴCy��/ڙ���x�}r)����ͬ��.��M1�b�L��9R]��#�P�S~?��~�S�h(������s��Ig99��.��"1�3#���'�2���kfɱb�H����#��hW�<���W�U�Ȇ�PhȔi�-�YZǖ���]�_�y����:����d��Q�˔s���X�Y?_-�����[�,3�"���e4�, S�/N��/3R��o@GHċ��h'�{�lQp���b��nB�{S)@�`Id�!kH�iH�i��!�.�@aK��-�&�w#�@��R���ʽ��C�����{�9�{�S%�*����Z׈�nV2�WN������)q�tJ�r�� >قZJ�q�s^W�a�B$�lt|����j+������Q�^Ы�L.��O�[���'�Q{M�E���.sy�9v�����m
�6�����"�^����} &���b�Ě4B<��U����Q8�0;~A�mP�D?��F�O�S�`�A��6�QE4��A%g��?	�M��:ס�ͦ�_��֤��c<�S���Q�eEp!eH��5�Aq,�/��b.ō�9b�.ɜ��~SGvO߯׈Ǳ�_�pTj[��5��w|kb�:P¶���5�&5w��ύ���p�啦�%����;�h���Ϝ��a��g��	�W�Z����d��]�7�ma���u[)7�/P�E�&e ��]i�D�P�t�J����_�:���^�qi���*p]�m���~��Q�m�{���V'�.Â���$`��,O�S4�ԋ�Z��[(�X۞�^]����8���f�N��ȃ��]�O�~I�H#6ae��)��X�P� S��~6�Dc���	��hV'(��n�����F�|���[�f�4���������I<.M���Xs��/̄ښ2��ͭ��/�5��˳}+�{BI,��JF�Xv��� �'�v#���fA�!G�R	��"O��p�|�k���&�P��ƚX��%�!�P�pv�/GO�qLZ�D"��xO'�C	#K�
�h!"���gw�z���KD�;\��-����}��P�&�u��p{�q�b��'�Y�I�~n����s�������q8����垜����4��ק�O5? t��0+�V�`<o	&�4��`彜"+��h:��K�{�s��]�0-^m5�k<�W;�2��S���Hۧq�>��F3���Y7�k��>*�!PٗC�1���"_yݝ%}��V�����6κ����15��l6��c�pEEU��:��{C�k@��#\�W+yjk� h�,+Dz���D��0WdY��Wn�l'��^K�jd����a1�ln�n+:	j�'��x�_/˻z1��x��b����,Ӑ.d84�N��P�GD�y�!��X�	h'��z.u�%�B���FS���h�7���l���~�*�}�C�t{���6�Y�o�s�6���i����-;�+\�H�s+��L��"�Ѽ��;���4����N*�h��̉s"p�I�;�g���4Z����}-c��������W#ү%����+�;|?���Gރ"�	��9g��w�j #���T(��̉�_R���/�L�N���f�0����r�˳��s��܄�ܶ!�ɯ����
m	(Mjd}��KW��(�9;xZ@ٽ�ĉp�0M@+r���:5���N宴�̧c�Ua�*ǊW�҉~����L8P�NQ��Mv*�Y�#xMW�u�n��pX^�f����$�� s�'��y@C;谹 �F������p�w/Ebc��?��1�?W�?~ሪ�ş��cͽ�>��$����~���?�]*��ȋZ#�3����K?��~z��0��`ɯ���7�NY��7�g��֒�)|��	�4�v�P�ɽ�YnXS�KJ��$0;��;w���qx��j&Xk�
:ˬ穿��I'`�Ǩ��K��Q�O���Q��\}Du���D�y�rg�k�O#/A\��I6/�+z�H����H�兴MW���8�Q��Иnr�Kjh��#�<Ī�EG�A}�>�������:S@KV�:z��-;�zPz�y�%�\�+!6j�ޘ�7n�l�	�@�g�Re�׎��>��l�nٙt�m��!�WN����p-�Z.T�� ��C\\�N��\b�	�L���m�g���g�F5KI��$�'�}��P�έ��P�����c½��|6("��Y��M|�������� �3��f�2y���k���O�xکH,i����G�/�PS���s�3w��{����S�����9���V=�V�f��p3�F�^huYT�Rƚ�q�؋g�bЭˈ%M>V����5�������k}fp�C��i�T/-Q�$��_r�x��ӂ]�Μ
2�\̗+ʤ��m���c���"��WtbҾш18_��Q�hL��+f�^p΀�B}�ǭ�Ő0�NJ8z׋����?�D,���懞Σ�;^�P���{$�{�����D=Gu���Y��ʹ�?�Q�6��D�ʹ�6e+�.۶�1x����g���#׾��P>K�@�����t�%�rx�^DQ��TZ��S�E��E�AgMP�2�Z�G��U��-� ��AZ��y���+�Ӑ�P�U��o�[�Pʴ��j&����_�׭-�e��{�Aa�+��6 ۰�
�Tf�����,[������M-77nM%�.�y�?Mre�>���z��W�P��FҌ�
�h���Ԛd-h��l�R�>'vQ+���#ْA��?&<�[۠�/���m/Usm�7/:.��W�Cɷ���[*m��\B�
��D��;; q9޳{]�V���?mg��v���Bq:�w�N�?�#��C��+����9�^����6�%8`�y�+��GyAʋ륵��,:�zyHn�I��༩Y�S*t`���XM<�Z�ũV�T�>���<���&":oV�T�_����[�&�sb�Յ�����l*�XD2uܼL�S�b��q2�JlW��E������:kE Q�fkks��%�cb��
��P�!�0��Az9Tu�8 ;]�,h�R�y��7��ss֐���ԎiOI �D��Nb놕5��䨈e�h�|����j��sfYK��j��U��*z�`]�K`�vû�om-��ϲ���$s��s���]�P�����ɧ!�|�2(�~6�"�P����\u��l�}8���j[�өU���e�2\�z3�p�\^�rV�����r������&�x���2�I o<���zrrǠ$�̽�s�$�q� ��W���>�Ҋ��o��3�c#ë�2FoJ�℻}�#�#�� ��N�H_��CLp��� ���������͎g_���m���6������ ���Z�����L�}�>/	@�;]�\_.���cx��"������(���ЛO���ڙ�����/=1�k�2ڮ�jߍ��� &;]�i��4Ve��a���Y~��LqSIdm"�D��$���x��1�rA- �$l��Ln����4�,�;���+:'��o���g� �}H���s����b��̬��YU	� q�^��\*Ȭ��;�-�RS#����4��Tr]q
�q@3��ox��Ėݥ1?sY�Z.�<���&'�T?.�c�D���	C�~ʙ��S�dr��� s�ht.P�8�2Q� ϋ4� iw����5�NqԻ�
}5�r���:ٯ�#1�՚�/��\q�n���O?MaXf���4#�<���c�:u��i���EĳZS�؜]~�u�MOF�E�����3�U��
-�c0�iz7LM��0���,R��	 ��ΫӆI�==�6�~�`��G�Y���w:��.N�b?VB�遲���Lm� ������7���mW���e��y���#W�\�Ou�_����F��OV((�5�J=�d8�ъ��
 �6���	<WYi¨�`l���������
~�Gh��9ж,
�
�\�5��C�X\M�E�كf3� ����:��C�`R�g9w�2�����x��{�=Jz�w�m�f[ܹ�>�¹r$v��I���a��ӱJ�TR��o_�:�L}�3�Ȟ��ۯ��ET��N���
�~��\�-?�lP���!:�A����Z#����!��o�"�=�쉣�%h?��a�@(��8+f��X�'��}m@Q���R��W�e���Igh�M�D�@{zA������!/w���-V1_ ;J}DP�B(���B#f $���Fo!aR��|Y���;F� �[_�.|�!���7s7��|�z�g*N��4{����^J&��B�#o����z�$W��J�)�����kM�LeT� ;�gL�0������?1;�%o������o
�/��d}*7��7������G � T�d�<E�>��V��z�`�K�9�� N_N(��%�s��c._���(JJ'�6��j!��?��+�1�'&���,��3m�2թ]� �	����A �`"�xx�0�� 8O�D�6KW��2��m����0��bM�aYN��C�4ntLl���r��VW��%rl���ySa'Y�IH�KǙm�?�e���y�
ղ,,~i�r˭>����5�RM���y�oi@�����l@TE�r������ߔ3���α�`�Ⱦ�/�4G�|���vr�s��2�;����v��iT4x�ܑA�J�R����7�{Ѵ�u�5�OK`5f���|����nPt�}Y%��R;s<*��u\/��V*�k�ǭ�6!��V��Qb�O64��INg\%�`��,���x���H	���U��)����_̰,"�u����>^�����g�1�Du�w
��f�m��r1���?W��ў:�?5�% ���_������5 X��#A����_�-z�}��;����ȵ+^�h�����Ee�$&�O��M�B'S��K�+)�,��3T�G�2��Q��놨I���@d8�U��w�m����=��L�0$�T��ht���7���4��$pB��|N�'7w����Je�������ϊO3�0kH��ɑ���s�Ҋz,隈�ͷP����[g����Н\
�U���xA&D�Cu�顐;��_��z@fY-�0��V�8� .��I)��TL���-��ÿ ��o��Z���S�T�.<�����`�I�5�trG{�� >[���������XC��Wg8L��Y1��3P)e@f	��;��XJH%���
 ����4?x����`��	�ͦ��,���}����}7�gU�6l���/�r�]���R��.�2�����bO�������4ꣅ�6� ����t;�BtCD�;�c,8���Z���dR}PxkG`�M�������_�͡����Q3/a5�k���٨A�]�,�)"`hn�ǟ8!��ZB��N�@=�,,rt��h��x=�p��D#Z州ׁ�?-��� q>����:%k@��\Q�=�0�0MĴ<Fx�88�ի�[��E`e������K��ӿC(��ĨE�����ԡ����]ČJV��y��q��_�>�G��n����^�6y��MĜL8i'��)=��Lp�ֹ@e�WK=�����\���r�za�l餉S�B"G[	��"��� i÷���B��)�=&�~mG��z�Εqb��y
J��`n��	�*kS�}$����:�w9�F�����6�����-��"T�>�}vd,���{������m��8h�e �C(_�GI�R�y�r�D�j��ϧ1�������	Ù�1*(Wx|� �W�~���csA���g�l�"�T(�X��ϧ�ֹLzu�iZO�5�S�:�,�lFV���K��}+�޿�Ӏ�/nQ��`�)b�_Mb9����1�B��WrD|�C罷U#��$BD�����e�v��V��P��kܺ�?0I)��ߎ���gH�_c(=�==q�Y��:=����|��w�%'US�S�fR���󉍌���0��a��u��5�oIߴ���$6Xi���� ���!s��X�������Q�d��G�� �cz�G��M/���s~_�g$�H ��2���Z��.B;򈓀��/d�jBl���T�e��Y�sz�8���	j�σc���E���6�˗��̿Pe�� ��4ַ_���n�qH!�N�Fqc�=��v>���
p���f��JC줉"��`$@G^��H�s�W��F��Җ�ʭ֧C$#�ZЀ�Y��DΟ�L����N���G肫��q�2e
�>���*�}�1��� �.��I4��F;�#O�������m�`��ҫ^X9��r{d�B &�I�`�V�Dvb��W z�f򲟍D؄��$�i*���O{m���{'9?!y^&G�KܜA2�Ɖ?�.���k��jsh4�o�ڸ�4d?�#"J}ŦHL�oĎ5(E�#����6�i�A#��7��_:~���Dʵ}�Y��L'���(�5U@J��W,s���h���ׄ�3a����x��m��\Y��ϚY+b5�hXr�	<e|
=/¦*���O��ޣv޼��
��q��4d�S�M?Xh�y6�\�`��(���"�E���{��;���q�-Y��=Z~�g=���7��l������0���YZh��޲��J�>{�"	�Z	p^�2��'D��3�?6���x�^�m!�|�愴'#<�L`��=�!�*�l�4�F>��;(��P7�We~�f�+ƨ������g,�A@睞���ܓ��U������՘�A'��_p4�b�͒d�G+Q�x󑇹���v1	�FyF�^��$|� �s���>cAU����ٹQV��A���� ��L�>�{�PH��T-�]��|2O�^:�-vRF�Ƚ��T\����e}*�E �|I�\�JFϵ�����hE���qm��$ޑH�.m�H�z�g5#�Z-裉�6��o�����q���#+�#󳻐�Ȩ v�N�|zp_](/����B��YU� ��}"D��]�W��m�AtW�rp�)�V��s��w�>H���L��t}�c��l��Im�"��{�1mZ�J�
�l��L�+��28�zm�`��_U�yV�_��*������q����bKsی�
����M�G��?J��@i@��,��c��r?�]�<�?��A��c���v:���ǔ��[�Y�lw8�ɯd��~p|�\�2�/T���4əiWYCf�jen�}�^o���<I�؄��sM� )���g~v&��{bn�b��jgrϛb� ���	�Mҩ����0"e�K�L�`P�)��c�a�GF����b%���'-�2v'`Q�XW��6�E@�	��[�[z#;����X����VaB8}��'.�!��9T�@H�aX�n��s�#*d�uO�ǇӲX�4��ѧe�҈�8X+�o��K��Pt����S����͗�ץpGl������Bح6��i9������0�Y�z��y6��JD�$�օ�����S&��hG9=Qi�aD����6��L(��o��˷�D�����p�a�0��U�"�l*�z��ӱFt��w�N��x, c�{{�L�����Z�ީ �w�{�K�F��D<N�E_3b)hW~��;���?��[RIi��T"ɪ����v%���.�1!���Hw�7'P���˝�B������z�����c���Ihvw|����g� �+��,�~����6�`-�y����ֲ@��������[k�j/��K�)۞�w���b���fb�@�����BY��E0v��ܢȐȒĊ���I���Z����Kn�;nԤc�)��$��0��e_����J8�E٣OE�-��Sm9w����o�<*q��]��"]Wّ�+�_�	ϼY��^`�[�=J�;�^��y� �)��-�qi&	���ҞKj�L�E2�x��c��Q��?!LiE��Y>�%~��Zŵ�]0n�v!\�5��R�����ds)X�^����)�:�)��ٜ��6�]�c:�u��c�̌3�o$�@�m�v��S�8�{��w�D���]��Տ���yc~_�e����s���M��XT �9����
~�d�U4-�|;�w��M&�M-х�׾�����:��e	Q���A�p��pK��om�[�s K���'Y �]��ui�m��te%������^��ypP�/�E6b�](���>(�p��?Ʊm���K�1'��f�``��J����G��V,c�U�N�/�P�}�Lj���~������`������~v!#o���PdD��TX��+&QYl���9sh��7���K]s�� ~Ϋ ��h�c�&�b�ތ��^�����8�̫ex�Ҥ91H%]tJ�&�� cV�for����7ô��`�hP����*��=�*B8�N�������p|-����fnb���G�@o9����,&\��<CH��O�Z��V��q����j%-u�R�������4޲��zM�yO"_N�2���f������D�^3� U��m�Lw����of̱�S���t�i��~?�H�'B�t���޻UdY��[}PA�:�U�W��쐍6�)��-\6W$u*9`q�A_�`�_�v��.?sj������p��M���偮u2��:�%9�\�[=ʅ�ث��W-�2{I��Tˌ.\5�j��?�����|H�S= n�Z���U۝M�,H���aJ.AI.p�ḧ́��J�
X���=7��9��a��j-��7\�Jo;�_Id��<�I����o5��,��f��>R3�E�y��U�|a �,�{�E׈�߭��Dr��9�p����@+(0l����E�s�� �䊽 a��fT�;{s��>�Qp������$���}r��.s׫��:&�<�{�`ā�dOy�y�}�cd6r�n+��f�������q��eCg�&�����S��;�D�� c �T�/������,h�lY/tJ�p�� 1F64�dߥ>�d�AY*|&���S ��� MN��0J��KmY�51�qc��f�Y4?,��ޡ��-��Vķ'e�JLsc/ds��.{�*�����\���SY1�����D�)e<2O��%�$���8�J��j*��J׀6��������ǭl5\I�;圜���1Hv�==T����T�v�H�9v��0�Ifw��!S��g/��6�O{@J� %=`��K>'C��E�C���͵�s��u�>څ|c���2�f���]��=��l@����$Ԣ�_#�|N�!ó�t�u��ZB�?���ս��1��v�����,=�ԉy��ȿ�p�kb&N�2Z�o���D��_;g&ဳc8�[{ʓ��!C��]��of��K+�Y:�і4�f�������0��	+��l�霂>]��.4	=�7ח�K��tA^x@�Z���=�b��SP���%�eA���
��Б�MfƩc�*��~�5��k�&/�d6ťP����q����I�|_\Zf>ZzVV����(�<le~!A1
y�u0{eq���d^�B2�r4��$Q�%
�o��f!��� 2$A��g�aY�<3�8O���V|�Z�̬�ڹ�%����^��5�f�9�#cl���ܭ�{��H3�|�,�'/��^��/1��>���f��Q�Ȧ�[G�u�],�8]73��^l�b�QG昦� >����:A1Qa�UՑ��m3ҵ�^݌�B��ٶ��WZ�üFt΂��OA�= ?`��b�����f݄�@��2��-w�H��Q�%{2��	�i������G���b���Y��p���X�K��W�xn�`��r��fR�D_�%=u�c�Iz�, �d����VK�a�y�R24e�g({�fS%��k��[�	��ں���t�X$u.-ݝ88��g K���S��<$���f�oM�e'�3e��M����Z���6�&CQ���(��j��.�p7i�΃�$�.gF��)�6C��p�ĞX��l����[���a?l���|AP���Lɰ�gf&�����$^��'m�M�[o�)ΕRhBi�������� 䥝U:�˕NS�"��p��'e�,<���C=kr6�t��AC���9�8t��� ��
N_�X���]�J���#S�t��}�"�,�S��yq86[��(�"[J-���Q��20HN�Y����QGV�=!��\2g�`[�"�!]  �n��]��R�&-O��Z���y��n��x��:�A3��B�~���ٕ�JlD2�X��+�'�>��X�:����oz}�	�p]�{�G�K�0�xu���fp�ڲd�]+� ���Hx��n9=ȭ�[ ���C�IzS�.˜G�M��R$�ǥ�.�cP��f� ����hv����{D+�t<�#QYcG̯�W�f��ٷK�8��xA�	"���Z=`��嫧,��_����`P���.�S��0:j�3L�8����@���̀�غ���B�G�����ME�?ga����+0R��&���.J(�w:��M�١՞+�[q��ெR&�I�03W�H(]�/��ݴ�!��N�$���	7�j�,����G�m=�?����WA�$D��^�]��R�u�Vm��Hu�k.��
�UیE��CwB=e˘��"eʕ��]���I�S�e���I�R����zb�[�!�Х0�ug�&ԝ�_���3�`���'�XN�P��/vD����/s�V�+�#��a[�����_���21o7D*N9P��#V�R�@�e�ի�|�@��Mr����fiu�+�l[Q�,Y��.E��7���M��=�'@��\Q�Y��~��~cC����f�7=����Doi�9���NRwO��S���X���R�_Fg!Px�z=����'w���&�_Q��4�m�I��U��Q=�(qƼ����㙸F<� ������t�|�|;�aB#sl4��ɓo�}���_w�w�aZ��MCY̢k�	d���`��F�7�wcGKW����̂��6��1`Q�r�8�w	�Wf:�����#_�K�ۈze��@� %�������b�����^3.�*�����}Ԇ+P� 8���5|�fKIg/����~�c�:ʧ�Q����ŗ�6�����f���8]9A�ϯ��i{����MP����o����	�i+��yeE�N�}<Ŧ/@p^8lP�I'��OS��lN+H��j��'|{~"C�Z�	�ۭ�uU�P�w�܀����(\'�W�t�����������j�{1�E%~]�bΑ{j���5}M���*M���#yg��WN�rُ}V21�W�����bm� O�iE6*�4d|2���-�Ezg�v:��P'{��PF�N�_ H�$������Ճ
|h�f�-T3��Z��g/dkq�Z��!��x���ճ���!�(/���\��=#���f��+r�a�^u�<(,I"ZҧZ����:�= �$ϴ�J�}J��R-�y��pB�DY�5y���}��M�NV�h�>�P�r�J�� Ƥ��=rV����P q���@�a>�)I[�z,��u|��mx�h4)~	YokCE�_�ք��Q��	3p	�`@��w�)��������Z`�}xOW&�����k�s#��L	u}.�/#�)��k���"�j>|����+z�8h#�(8ld>���$ɶ�ҋ�{r��Ftqz�o#�)�4�hO�_i�(y|��c�W��h�m�"F�WZ>!Ű�#�ͩ6���B�/ą�ԩu~�=Z�k�m��)ysoxz��N
�@�^��pZ��y󁬌$>Dx����zSI�63�)J���P�s_����x]���$FsEKц��@�ɞ㓱�i&�є�A�i^[ʳX��N'�:U���M���K@%P���Ɍ�3��1z��
@��}� C���n�Y�~Y�6ˢ:J�t����DHݫƺI�^��F�)��k9@��/�ϣ��rNB�Y�5T�h��9
b��]� �Sp�ͩkh���`7L<5%O�\�_Qw�7���4�=����'�$脼�(+����v:�s;�?��v:�RL��핪9�]{\l5|U��du�I�RR��+S�=�%�w���PgӨ��ܹ����fy�Px��td��]mC�zߦpA����f�2�%��	f�߆v��Lw�Z�ָ���1c����w��l�������Ym�\K�Y`��~�����.�Pj0rq��� ɖe�|�γBËx���D�D�-^�bm�V0ض�i���S����.��Uc�h8�(�a�T��UW�A��Y�R�q�������?��eȵ�	f���������6�_�������?ri�v�����)],φ��y��\:ᫌ��g��>�Nu�<�hU��"�LE�Y��d_T�k��������Bd�f� -�@6� oh�Lֲ���l%��(j	2NOxv�	���ϥ;5d�ZºP���|��ѩ�"."z��Q^qA_K�o�>��ɈX4v=�۵�H��}��߸~�wI
P�r3^���h۠���"��Xh�z@޿�G2�i��Y�F�ٱ�GNV�ʕ��	�$IA���X�9-�X�S�n�^m	h�~����}J�*7�3ԯ:L��0��w�[�@Ri�AEg4湃�����R��:�N��������)>�X�yҧC��S1@��޵���'eE�AU�[|���}�b3j��)�|��'�be�k�&�*��Dq��I��o5-M��['e���إ�U��\G�7�a��z�+�C�K�{�y�8�.�쟷r�S0$.�L�R�!�=r���t����Y�("d�Iڇ�Et��=Z��rN�#4� {Y>�L���?'��z	���S�=<A�e�f�a�>bk���<�y$ ,�ҀdL��|�}BDL�xm�0�8j+���w�n[bn����Ҏ�P��L>�18n�4���vڭ f1�o�휗����Dc���\_jnﬣӅ}�rZ�ym�2� ="OY��>�[��>�%˻���87
�8ޢ&�s� ��,W�9��!t�:��S�_7:H���n%>���=�����~f�����[ �v�:ڬ܏�6����0]��IE�����w�l��*é����7��.9އz��O�S���k<�I �e���C?��n���r��Xv
#ҡ��)�jj㞓�`5p��?�C��M��[b'�&�"ة�@A�z�:)�[�>�K�^�T
�Q�ş�p�uO�GY����:��)-(����Hy��t�7�����I
I�]�B_�e5����������nU�� Tܞ<�uZT˄����۔������K�4�ك���_a�cn�{'d�5G���!�z:�z�;�a��n�e$�Bm�����@�(��.�Lk�cg�K��5��:��������%��� Õ�A��u�rиM,˃#=Ӟ�i�@;��+�s�#NS#aP̼$ҭ��-�Byl:����0���_Ű��)ǧ睂X�pwU*Uln��-�P	���%U(��~պy��%���8\_��=|�Xk��<��=T
�)[�uSU�� c�;�;C'>J��G�`�,L8�1��j���@��*��eLۋ:nk#�8:}[�Z;W����>�c�~|ߺQ�`����Z��qSA�}����]��>��n5�A�'�(��e����2��	���/���p�-zN�)$BjP����&�J�~Oc�ғK��U�	N�>C���翉.�Q�f�bU"�w�����-���u�]�7MG:�G����n'nrg}*6=L�[ǲ�xe� ����Q��ile:�$�w]l��:~�k��*��l��f K�m ���� w�(#��5L&]�4����r(P� �R�xG
�3�:� 7�W�E�8ۀOj �fz��k�H��!�eIs#���|7����v~-�B���ɧ_�6�t��7~�Z4�E̽䩂}jۙ�q�V�+	���'����c�k�<�M�ňځ�t,��<"�gI ��3�b���-���++F*��y2����S9�@H�b�6L]_Ol��"-\��7����]��
���-�[�(�#�
~���'��7�>�U���F���1�$����N����c�)c�T��^QH��NmG6%���	>����%�3�fh����*�`6@�3��<bi�Ѩ�y`g�X���3сlB�f��6�˕�#�n�>#Jz?I�����
���?<:�
��{�ss�K!��Z�*�XA1�yRs}�M^C#�kO���F2��*]9�G�d�ϼ��9V1Z� SMt�"�9���[]�w�%@B�i��o��y�(�I^��v���*�������
�h�T\�!kJ�t�� ��H�ġ?֔��t��D�v�qW�W�27kH`oM�m6��"v���<?-�!��X�|�|�P5���a�4�l����7b�u�|�y������̈́.���2O|���/�?y3k�q'/�ܒۏ�L�0��R��\����i��n��7����H�����>X���ʢ^d��٣���!�R'X߱���3�u1b� �/��ja��@e��q"�
wK��������#9�(�@��tr�t+�P0d���=/<>gK˓��
�Ŋ�����98�Am3%��|{q7�6�D
�������2]�����Mj�0,G�-�'�0m�τ2|8��&��N#������������#��H�*���*��S��.�%I"�2��F����S~��h�\�.�+�@�����G�4K7�����&�@؆Q[O��.��=��l���9���J��g�a�K�)y}�g��KX�?/�k6 	�_s�=�JKc��'饽�F�?�U�5��юξW��}%��>�]��T��������sʤ~I:}��O��<i�^��W�{0z�>�_$q�a`�6ѥ��wu�O]�
���bfu7n����$�`%���㒿��"?��	�W���I�&9V����t�7EW�8�w*`\Cs�A���2��UۻzDX���H`�}���/=GU��웙�a��L��0ك�´�����!p��Ϲ��%pH<���#Ͱ_�w�F�C��M�.S?����hD:W�ץ�Ć���2�x'A���Q�<�:+"��v�-��.I�$ `q�c��J�։�-��^���o}6��W�>`�Ԅp�~Dã�We�Bz���xĞ8�흡%��4�'�#}j�S|r�c�=�]j���A=W�/>��:�*;n9�ݝ��4�m�
�H���(]�W��P�����3ɿ�/�#Uʴ�xTO�:m��oMүC\���ĳ���}<3Y�F^J¤IE"_[�QL��°�S���Gc����A��$0�@�pn:FtĆ�T%�-9��D��bNx�.�����H֔ �K���7��P2���3m�E��F�+ؿ��Ew�=�Y+ �c�����2j����l��*Bai�8$kNVz-��O���|�\��w�=`���X����z����l`S�ws�3��M'�p��O�b����~�!��`�t�MY��<ɋ�(l���h�L�+!��L��?;��s�kh�YH¢=�����B�f�I�U�H_`i��[(�;<�����R/k~��ڃ%,�	ш��,��;��`JzۜB��2����&|���c�G�>~<�CMT�.7�����#���`8�N!�gǬ6��8��s�PBmS��\G�g�c�Հ��P&�f��s�O	�DԨ8H�|���(-���%@1��m3E�H�S��C6���5�&��.�X��Q���:g� _��!��.�"P���k��'�%���#-�戞nh�T�
���q-��;��NҒ{�����J�(t�������?����v)f�\�qT`fS�u�O�����Y0`���)�Xr~�	����y6r'����l��=�k�]V�|�+�1���˶4��:wz�����G%��Ѻ��4�EZ}9m7B��cZ${�d���k�@uE�Z�����h֪�k�`��0��G�d{�H!�EQ�Ot*��r=�q��˼�'&Ho�,��_e�ެ`k�)�z�O6�Z�~In�ƇLr���d��cG�n�ʟ�!�
�]���hǙ��������m��3	�ȩCZ��j�yۻ.�*����LbQZi��喓w��!�T����MË��_�2g����Tӌ6��~�2aD�8�����0t�{DK�X�����Ӵ��M��k�L&��j$G&I��
�g���b�~�hb����s9��=MC<Jt��Q~��73>�x�]�%�N
���m�#TeQx��	9�6P�}��u�egc�O�4��>���$�J�M�H`p
�Tw!����*smm�p`��~E�.<Ҡ!��S]f����c�ց��������k�p, w<C;׳�Ս��N\/k1���KA[~n4�>���>�!1 ��<�o����l�����h�'c�x\��Y'��^�}Z��Qn��g�(6Bn�J"$���[S.�g�[3��ø�
u5OOS�7��h���Wb9�\�hl��i�A\S���;M���aI���H�s*����֌L��"lU�+.{�ա��zŐ��geU�/����l�Q�������$�,����S�kà��h�yh�Q�13O��V���=���S���b�K����ۇ���[ �J11]��l�=��2������N?�6���\���������@��w9&Pr�)���d�F�,o��Ǭ/�#u��(��Fv�S�q�u����˪��=��w�oXi&U٧:�l��R�hU�e��mV⁮B�e�sNZ�������Cf�Z�1�U!;p!�Z<С�s`jVa	_ZP�+�9?!V��}P0y+nAT������*���p�)�Β�������l0Ua���g)�,�FH�Ԟl�Y�����q��;�ҧ����A�X�OA1.挰�keRl�ć��o��kt���Ǎ��m�L��� $uF��m|�X�AՑ�`����F�̊�R ,o'�zR��B�_���WM�^� ��Y��&���$����Kc�xASt��˺����D��$���V�Sƫc)��v%���Y����T�;gE�����+<�������p�Ji�J�S&�E�C��K$J{y�+�Ζa(I��V���|�y�/4@�nGO��u��I�>Y���"΀ �E�Emy�t��绪�
�z����q���3��Y�sTfIzߵѥB�z�v]�u�Nk_��37 �u	��)���<�����Hk�|wZ8�'a���o�Ѱ0�{ַ[q��U7�{��ۅ������y�J��N�m���E/n�����Y���r�We���8��z�o�4���<I$$���w�*P�������9V��k�j�6�d�Q�zW�VB�������{�$?7�cŁOҎ����,�Y(��0{i��_Hv֖��w_�]��* 83���Eb�u a�7��;(ʖ�����R��>��0���'[��W!���.lHU���>o��k'�"οH���>bA��4 ����3t��Ŏ�}���j�%D1z#��!|�]��W�.�Y���e�Ñ�5B�����W?� ���Ő0&;�(��I.�A4G5�!r	����@�-�2a�je��
��r6�� \1S���q��z��s]n�M;�!:G=
���z��

w,�p�¼J�<�����R:�O��ͪ0�h�Cb)��͑"F�$���s]��*�d���VuBwDx�q\�д}'�C��Lc���cbF�؈&�%����p����=J��eW=�Y�XwR�^��<N���ʭ�J���6ÂY�Ij�<b����O���<:�,>��^�cE��G:{h�����Inv,@rI�0���B���+��.�t��.C	��j�4Qޯt��U��:�L)�ي��/'�yl\�H��"�?eNY���iç"�h��$6o��O��6| Y3�p:,8${��娫Z*�^Ѷ���;�����w�_�i�.xvǈ���~Z|��u���c��/��Ʀ�>"L6êgw��ũ��V���Ƥ�JOi�U���p�[��*5���v
�ﺩ���Zc���np|�SJ��ڍ00h5S���H�p�]�~@Zl>�IF`S(P+P�:M��\F���;e�R@5��I�)o.Ԕ�0�.0e�4W;��"��eft��U�0DmWT�?m.Aj˯�2�����\Iq��+���9[���iP2[q�x��]B�.6	m�<32?Ѻ�. y7���ApG''#%y��HK�nO��7�����&:�x�R���`�(�����;-j�݋r~�\O���1�V�ǿ@�oh�.�վ�����p�P���]� ;/�xu�7�dOS[ܭɂ�Y��R�!��v��9EXȀ�1��:%����y" �o$�nH <u���fu%���L/�}o9�yG�cLvc����X��X����]�I��z]C�vm���3k��0��D����z�ۈX��<�]''34��� ��� ˖A��U#
���,)���f��C�&�Mb�Z�m�b��M���-��H��=�������C喸hM��:ߔ9��咤�ب涉K��ݦ��Iǩ-�.ͨ@��f����!qkC�܉她`�K��-Ep��.?��z��$_{%LQ^���d;�L����^>q�ڎ�F�oN�9~�y,%a��RlƖNX-�������|�4�Dѐ�ص��L�t:/NJ�SJ�9�i����5]�df�B���-a�A�ȴo�����~���n��)/ �ݐ= �ޤ�Q۔�:e�|�K����.T�9H���'�
2r��,?�ȴ~h�'V� ���<9�Zs,�c�W��Y�
=�1S/�g�I��*�e�I���V� 5���kpj���2��5H��5��w�,�ߖ_�%�+��Y��p�aYxmdE����8���S�F����:s��P��%��&ܿ�� 43�tI�2�9��Ɗ{K@bi�cw ���*�|�f�`H��a<O.٧䨼��ޟ!�X%��<�R ӝ�`����mq}#g��N�AxJ���\ ��щ���:ޛ���$��$��]L��|٬@���,��׵F~�d�̨��_�\�a�)�Ã�[�,�t8��� _$ �)g��eT�<�ï=n*
GR��0a92m����}���:�U�8�H���� ���lY
���v����|�n1�Ѩ��y�����1  KM5���H�j���. ����+c��1V�z9�ښ�G�
|	�f�A5���4D��"X%��]^�x�����o?��˙;��О�L��<�Pr�wgڑZi��2Í,X����@.|�V�-��J�a@=����O����G��r���߇�@~"똷vt�j�{f��� "���Z��^3���l��.�'22�h;k���4�y��Qy��}|oJͤ�����rM�0;����x�S�>[{ҀJ\���p�%�p���KY�eW-|��� #T�:7:;ݯ3�� ZԜ`�r�������F��)ΜH��BvĖ�3�����|8��?I��I�<NJ���R���M1z;���N�?��vEϣRc�lҹsIVX��P����9�^~�g�7Uޕ�]i7R�R:��D�
�S�Y&Hю�s2��Y��w\�U�N� e�q�+�4�n�~n� �ܼgoҵH�z+T����ĵ"��ت�������BP"���q��� �:�Ϧ!^0�N1�Ce��y������z��P���z�Z�~�1y��L�L;+xa�	p��'��4	��"��A@�΍U�N��K����)�j�H�d	�,-ς���`w�܃�mM,�٨ Th��¸uI�	'��r��5�X&g��7����|�*�&+Ds,�,�PU��9�Aw��O6w�~�����Õxs�"h�g�R"��n��C�|��mn_�� �u$k�/c>Yǻ����k�c�Xŭ��>*[9KFiQ��nu��M��i���wf�1�<�e%�5��É��cMt9AMe�DT	.!����1,��pO9�|��?'�Nw����­���%5�m,2S݄�d�!��L�yC����+�x�.��pU��券�Ԥ좚�n�+�z��B�
��Sv�˛k���ivV�ӍE�8�/��)8(US��_SW�Z��V�u��8��H���<��P�.�~��M|L�g����c���ky�F,d|���������]b����0͖Oh��L0�T뻔�>����ĵ��H�p4[7b.���@EUHY��h
��I��j��DMÚ�����&�N��,��yJ�����{長9�#~�<���h$D��#��1�����W�֮�"m>��3��*�W�L�x-�M��Ť�����V}�������+��X�)�f�u�G�����Vn��!"�&�k-Y;:��l�C���z�B�E�C��4za�H;-$G�d��ұ�/�rWo=�pT��R�A���oa����d��\�B.:��l�˗��N~����E0��X2�U���GR��:3�Y�U�-7��wa_�Ѝ�S�ɽ�c�  ���Bi �Ly��x�f@��̶�r�`G��B?��X�'W�4��"6�����Ps���-B6��l��BJ6N������9�1��w�`�ց��%�)�lK��j�*�m��d����i����ix�,�b�)2m��i�7
7���G�I�V���NLg���&�P����^{���6'��z���1���:�8G_�����s �
9
���${�S@ڤ�,��73������8R��W���G.�$uo��~���5w�G�&a|�<&���p[�a�ڿ�0T��%m�_��@�ğ��SA"!�,���%��z�_.B���`�ۥq���ۣ>���cd��]��9�bR{G�!��u�函�ӆ8��Q��m��c�I��'\U�M�v��'���q� �eN�Ԓi�x�zky�%6�_,�F_a�>�i�АdN�"�C?B�S��=]o����ܕ�%o�����suܚ���u�B�殏-:A\~��t�W��N�@�:��Λ7�i�B�{�U��C�/�ّ0�]��֫i=�"4����Y�-�ef�C��K���I�3+����/��G�S���p��y�'���xD��;�/yϙ��8l��o��c 1���Ҵ��+���jb��-b�;��2�Asǿ�`�~2�6Z�^b����^��0��'K�fՓ���Cq'�_�rt�#����2��-�t/�� �q���\j�(�X����'F���.����T3( �5T|c�G�Ci���:�v;�ڠ]�U&,x��W��Xf�F�m/4m��YyO�^�5�7��7k<�5��0���>Cp��| ǣ9-̵<?!�>�[�9;�qP�o�0龵��<�:�5�B���H����mY%j%�u��w����ڱ��"�,�Umι���`R5	���@g%Q�9��H �a���>u�&����.�!�s(ǐ�x1He���Y��oO A�`�T1�r��u��úEi���A,2�M�EÁ�d�
���|G��e�<�Mw��Ξ6r��^0"�b��L5TeT�
�Y�[�+�|
�Ö��7��)Kj�6�|	 =Z�l�$Puh�����ȕD�9kl _67,�g��/�}$n�~�k�@omf����#���ȗ�=k���� ���i��%��3aq �c� kD+ZR%�q����<��8�D�ӵ
i�ǁe)�3�K���ZK~��ٯ;�?n�(N�?���P���B:D?�\Lg�
�����gn(�k��[�0�q�h������E:D�)�Lz���PKD��0BA���d��HꑶY�K�x�`�i"A�"0>Y9d��e�{���x#�`�J�J����
ǰ�ݒ�`";+�-̈́���$�$��5f���xE�4�:���;�CU�P�\T���<Cu�{��خT$��]��7de/Ӯ�hD�e��
[�9�R�(	����υ9�i=�;BG�P,3��@����I��CU���9&��^����X�?Q��������ݪ1�NC�8A���9�J1ə� �� % ^s`���������袵m�>�ԙ^��,:��+6_)XL-+"6�O��`�p��X��J�p�x����f/�ky��~��=�8��|�2YTO�ď$[�=Se|��G��|Z��04���'�5��éc�3mW�
aGO(�
4����pAt���v�d�ш(���M�RT���Y�����]�.Y,$ �7�mH���A�s2����Z�O�O,������6C�\tP���7�'��V�J�N%�Bk�H8�m�6]�	��]�Γ��-7�!a��K�c?j4��quR��XBJ@��Y<ݴ�h�~Ԛ�)im��_��e��E�?���F��m_Ci�/�q	>gNp7�����U>mK��X�"�C��I��벳�BdWc*�R�Q��=4ӏ7'����=��0*\}��^�����P*��r���3���W(h\K-�5��XAN�z�}�B��)���j���|cl��K��o�*�!�3X��"�9��4�T?&�4�r,"g],��.��5�~^F�㕧�k�I��Sm���Lޮ� 3��O�-t=/��9��śIϙN��ݣՀ������0;��7��ߨ,6u8���D�̽��z�w���@�h��} Bt����� d`�����P&��l�dh^�ėnӉ�9�ʆ�d�u%�G������(8"%�9��]uQ��a���� d����Bb=�i2M�������Fni�kLR�o��M¤�#����~��0��!ʄXDM[O
O�;���9!6��ym�Mˏ�3}���6�a3A�/j�]��(�0���G��T7��l �KK�E�Ƴ�I��*�}5-u�.���6��47�E9�g�y�$/��꒢������.�O\-Ϫ�_I��/��W0����V\�3ey<�~A�F �q�^���܈����^�B����K�l��s�6/9���M�"�r�)#OK�2���gU0ϓH�������0�b�Q��L7]�tݣ)J�CS7\&�GĎ#Yx��N�1���^�r��F+�\ �H�rֈ>�W���e�u����?�L���HH��Y!S��|;�-rQf�Y1��@��m��'y/C�׏Rp���w� fd{ўp����*���~��K1�����+�r6���0�t���¼\�yF[�J�F���q���i�Q�*
������`��W;���1ԥ��l½���=�h�Wp\��M�Ǧ�J�e�CM�ϸ������E$��B9X��pU���g9�Z'�1!{'���U�{t�;�n��E�������TmO��4�Fir�Tܲ�=��s%2<&��|,Xi�uD�L�?�QFv�
��\�m&��l�#ّ�G�̈́i�d1|��N��Ptmyj>��U�ֈP^kA�#��t��V#lE�+5�HunZ��DPrzE� �l�CTk3�'�ޢK��T�4�sۨ�횓�����
�v���xV �=v4���	s�L�a���ƣna���f2��GF�+�`�8,1Ϩ���8�Z�j:�|�'�*�Ϛ��ɡ�8�S��Zq�j��byb�ױ�ƀ��ߞOn����WI���t��lX6�&sW�cW��	���ɸ�������B��𯫜�C�.���`�k��L��i�κ��:�{���@��Q��� ���2�y�߅��7A�V��1 y6��
H�/�&n��G��Z&��f���(����	s��!W	`@�\�Ub�k�[h@lHJ��v���j�V���Uƹ��T��҅�� ��Xe��$~З��i���rˏ8����?��DP��w8���,'WS�}]ßZM�Լ$��DዿW}�w5��5�n{�'�kMe�I(�Iv�'�<ELjG����������T�F���0=Ӯ���I9k��g\�Z�a���|�#~�G��;����c����DX헊���]�Ә,�ɛDR��|{�����Ы�`ؙ���P�8�/�Ս&v�a� ��ނ����v<x��č����y�~t�6Z(
��ؓw��*.�[��P��:�-��[��6h|��f�e����S��aBJ}�{/��1&+4E�`�q�d��(�����I%!��#��um]�at]�Ȟ��}�'�]���Ы���c}#�VH�νm\v!��C���Tӓ��~ �&P����)��JE�$�-�Y>��lP9]��:$qk����p��=
^�h0L�<�Hmj�R�� �Y9B��D�p�,)c2 ��:���@\2���o�ϐ92�N��p�[>�4��/���u*�I���&5��GS��W��;��>��ӡzB���4��G�'�AxD,�Qx޻��d�)��W�)�4L=�v�	NT���p��cn�y�3�Sa�h���]�(
H�����\w���耊�,�U췱�S�~�$��'福��a�%�|-}��)4��>,Q-���}߷�Nձï��Y$'4�TX�=�ŕc���{�-�`u ~T���9�s�#6nb`lߺ��$#�����tз�n}�	@b����� ���v
�z5Rr���m��@{.�qut9�Iw�Я��o���y���v���m.��Q4l3���	n��ӑ*������1af���4�}�t~l<�wIã�����2KЍ{bRdu*c$a:'�"�)08�kfw{�f0S �m��u[�T��!�Q&i��>v�Za����C�ZLC�9B3`�f�1��?�&�v��k6�"����҃T��m:��������]��{��Ո�!����H6�PB�:)ǜ��PP����+W5Fo�d/�-6����G)~O����2�BOOF׆h���E�ľN_�,���5�ƴ��������&llZ�C_U��)a�����z����/�mK�9D@@2��L��I�$�%��Y.F�5�W�!dZ)-B�c���t���PQ�mȇ�M�7)k/4��g�4��~�7݈�롯s�X����	-��0I���Ȏ�4dY�<���j*�м����KG5g& lX �%��c�� �`��7����p�S��nI�"Uy�̷ ͅ9_�{X���m�������M���+��x>vo��Qcd�M�\½a�r��2,�͍���bm�dL�Ayq����5I���Vx��}�g܈�P�4
6���Uٜ-a.J�K?K�5��TL;�ܪ�����sѸ$��.�7�m�&D�}��J��M�5�#�Ƶ�?����`��3���m��K_�l
��[��x3!,ǉSPGv�_9�4Az����2�p��e��ơ�Q֞ݢǆ�|�O{�������+*)e!�׈�ˉ�hF��°���#y���r+m��QY�b	�@���Y+u�-p�!qV�h�u��Xh@��E�,��7p<�Q��l#���i�|R�ɮl�����
�F�ҫ6_�2�İ@�Zʽ��lad���K@���쇁n��	:�y��/ZrD�!��%I�jI�(����e�#;��K0�j�{6��%g$c�&�L�.�A�0�&�ql �a�K>Z)G`��w	��O��?�����6i �=�?�n+��x�4
�GqV.R���5�Z��!*�V���?�����0�
�T'�2݉z����6�2�j��`�;h�θ����Ͱ�H1<෣y��! 2n�=h��/��w%��=���0�Y�|�1 ;"����S��9��4��oX��h�;7b��	byi3����4�Uݸ�!XXَ�1�[��٦~$�)�)lZ7(��%o^#<>�1MU,��o��'��h}��&k��U����`��:�x��LY<i|l,dM5��7�=��\��FGj�7����_#��v�G���������yW�&�,4"X��%��@�]<Q���6�{�����(���Y=�4oQ�z)�5��`�V	�%��.B�ԋ�/h{\��[�`v5\½6�[�~^g�$\�t=m�A?tY�Yf�e�Uײ5�M�EƈDǢۿ�̔�dbĠIϙLM����~>}:��(��T$���.�O/���d��,\�w�bϒc�H����\�����.��SHzw2��˹�a����2[/'����d\�k�/0*W�5��׫~S˞���m2��W��>6�a"\���@�46tsBW��:<B�~K�Ql���nXC�3���	�4F�����,��!�Ú���.��=�2�j�|��r�լ�yPI�p�7�(�I8Xw1oj�;��Z���x~��S�Ț�4O��������`@� .����0�];2���,!"I#�6z��̕�]�H��9�7���*֏c���d��¶3�hO"���߁=�`����2�FJ��;�d�C��C�M�%���3GR�xTM�Vk��Z%)�nJM��!��Rp�Ⴥ�v_�����0ݐ�]�zǒ$By&�~梽fOik�U�N�
��z�xH�4��s�n���`�I���������r�s�^���=Ih�В2� ������O �2w?z3J<�罢�h�(�c\�1@����J��k�{@*(+G�f���zr��,�e�H��Fu-e�����e���!�ܕt�� �*�&�$������=��Uc�z���7�U�.�FT���K�"�� %wAԤ��<+Q��s� r������M�Y��Z�eIuy��C��ڿ2z�r�ݡ�|���bz�U�q�zw�$y�e�����(U�X-'�H�%���MSܗd���C#Џ��{*(`t-���M��s{>��<��+%��b�4����9�2`}�>���# Rq'���Â휔���\b����e��J��Qcl�ҷ���`��Z��,�8��н�M�z��8!��aԿ	��9�z���f#a��GE�Z�Cl�-��Aܥ:��zX���Z�.ܣ7��,��Y	��ygK8oM%��}�w�Y�Ch�H����""�4oEo=\��{�9o��p{;X�D��E�I�,���1�w�(b����`-z\��*#u�[��$�����b�<e��B�y����?'g�ȟ�F�l�^�ȸ���JH�I��y�xyvnS�(�5�:��T��p8��L�ؤ�M=�n��r���Dp�y����e�a���ثfA��N��)|!�?C�OמX�aX�D�r���#����U���Kt�~���q��7�]d(�o���I�ݢ�рg�0�zaU��T�C��wOIEe�GKi
�^�d ��<tKI�]�<��{�����K��Y��J�b�7L3����66`����gOuƝ@t�"�/��/���U���1��?y�H�.�d�:�^����j	��,�!UK�`��̛JP���XH�)&��*E��� �:и�pZ$l�)��`p:,�B �I�2*��n���+�Y�(�b2Z���ƹcCĹ$P�w�?�g�	�B;�*�#[apV��
D���U��+ρod0�%�D-Fi[b�uՋT����^��f'5��fњQ%Wf��O��A�Sjީ��cH��)\>��}>^Sy���6�E^���C'd\L�}� [m\�B�f�՞�(����-����Θ ��sKtz�_FǑ�BMy׭��Y����'�[�hu8�8|<�ܾW"�ګs�4��9j|���Q�GQ���͙��LJ��Ϗ~d�^�$�E1����`Nu�P��S��	4���#��<AǛ�B"���Dig�v�=�O~�o�G�s��|���SJb�M��qH6��Xq��`��<Qv����̌�ILx#��}�>�C�tg�(�D�ʹ-�q�Ҵ���?���&�����]�~�KF�q@�o;[����na���tF^�y��t�}Բ�\��J�O4�qSD��8�.Z�m~¶�a	S�ǝ�7Uzn�e�KM�_\�n�4,�8����G&�r�����@h�}���:���L�D-�Q��H3�78�^a��Z�8"C��J�0�M����ƍL����J�R8��G=��-	3k��	*<@|6|ޛA%��%ϰ2R�[��"����~>o��ހs��%��m�j����. ��i;(܈�
W��r�&
?[�����o&�fH��.5��ZH�`YD�����H�E�F#���b�&Y|���3��2c��a`ּ$����1_n�R��=�����K�~�s]	X&��EE  �z,}� ��XjC�hܳ��>��B���V0*���n���+Ç��B�\g`���ѕ�Ա�=�����G��>��,j��ܟ��]a+d������p7��Z�6�<��eϲ�������qIH6���H�����-8���R�o?zDf�Mq>!�"��Em��g/L�7댧:�~�]�;�P�f�g�1v�4��|��*{`�`�옄�d�K`eğȒ��F�5�$�DB����v�u�o���L�J�?�T��Q)���4�p\K���7ĆR#EL4��ʓ���lA�,KG��)�g3���/!R/���ǂ��}�G����+N�����H�iMe+k�L3���3�����8U|�8�5&3�1K�G�~w����y}*a4����$�5W2~$���ξ�N�\Rr}�(qFG~3�07܋X�Y��v��9W�LEb��Yl��!v�e|�)�t5�����4�St�7�<@BF|���mP�"����� 3=�J��\�3�����_�y�-�SB�n��jE�p��}��� ��>HB����N����	t�:�v�f���&j���ҭ�7�L�c�ZM,���*�a[�/7I��Q����$3*�����I$*�[i&W кeՈ�%�0G������ޗ�M!�pՆOʍ��&IM4#�����6NYP{�tL�)%@�`��!| ��UhGf57e�1֤Hb�a�m<3���s����%8�}�, ���>��21�;-`�������⺥dCP-~�!?�69f~��4�9yr�׳K��l���e�~������x��h���ll)�-��<f¼RF�Yr]r��tx��9�C�Ṷ��������&���LGr�i�<mx9��U3f ��K��ֈ���OX �1���;�V���]j��O��E��+]�Jえ��Œ�L��g���Df�ӛ�MDgm롷 +է91� 5�ޞT��Q�!�����e�����W���B䁿����EdV���׵�DS�0�V(sg�P}�Y.�A���n����o��%�qC�i�����4ߏtj.�dK�\�:�%[{��~��1����z���W�?yΞ�uŏ�)ry�"��6��8��؜������1B��L^�{��3����g��
�멚|���ہ�c<jPa����������UWo�Ht���b���5�9s�A����P���!�� ��b�B6�����3�3Z�ˌ	\ӆ,;���Mr-�Ĥ�WOG�OF�c)�C�l9��<7�����.S��>�g.��ǧ+ͫ �ժN��`�Iz���'��'ߚ�s�D������@��v��dH�;1ҋ��g8e���Xy� ��r��h%�A6��$Zh��^�P�S���������L§[G�`�~��%v.��Y1��p	�-�uxý��i4����"�^U����=S�0r�����&��f��������r�J�î�K@,J1�D�->>��9 �cF�ep;�!�*|�7D����u������i��&�µ���b�����L��@z�2J�~#`%��1~.F���rRK��o��T�z�k�nJ#7��OO�e�H=�5�n�u�G�f�GB��9��E���_�z�B�V��[r.?D�CP�n z��֝��<�?�}*��&s�Zj2l��#���D�S�:��ND..>F5��!����9ƌ��R)�����)Ľ�K�g6�l��B,��JM��:rF���~>��-?p�Fw��*݇�Qg��τ���|�2B����i�2]o��9fl�[;d+N�ަ�d�Py���f�ꭐ��3�+O<�
�E�b�t�[��2l�?Q5$��#+���Q�C�ӯ�Ţ���}˵:�Y��D�?��dqh�9������:UP�v��a��D��!�� h�0��X=*
_�YK��/���A�o\�7dQ�ï<(d��J�I{�Ga�I�0��q:'t+~�m'�`���}�*��n}�����$�We0�Z���#�Ѓ/�XƅN,3RҴ�D�=�'{P:�*���L%$i'�Q}�<��&n�^sC�ҝ���.y wQP���}ʇi&�a��T����۵�Q���ћ?�gʸ�ҫ20����e��%������O�A�!#�U~ ���[b	�p��Oks����Uif����8�\́��z���j3i/���C��ՖtVI�U����Q�F�����!� ��i�P��|:��2N�)T��S����s���fd3�@Ŭ]�zI2�d���������ɹ{�jK�NQ����~T��z��B ���Iky�ߴ=p=���?E��&���	�ZS��շ����D�/�l����qA���1� �~����!hmOʐ�-I&����쁎0�����ZvVv�L��9���)���zyB��\�F^�v]P�]>��0�fSZ�YY�rZJ@�Ϣ^�Jg��?�;q]�ն��@��H�j�N��^��l��Ј�'v�V��D���^�y�l�Ƣ,��/���誥o��Xe�P��"J��O�98�"��d�r�x��(-����	����^w�ݑ��Jl\@��+*�1�l#O����[c~���J��Q�W1����^*_���r+��㟛���щ��{F�c��Am�m_�CJ�h��?�3y��6�C�N�	T��Z�֑m{���/�C��Α�
V��g����u�k�ŴΈUm>u�#yd�jOi�u��x<�;I7F����c���W��Q�� `�^BF���Z|���[p_���Q�����l�\Op1i��=���ex�����d;2(Q������8Z�>�����CA@���y�q��;�䇱�ʗ+Wl����䴠s���Y�
��:����>��/��'�Я�1J7o,%�tOw<��b����f��$�~�̫q^���}���P�E�O��=�[	�pǑ@� ���>�b~#$rE
*^p��qH��Vu��b{�.�B�����������>�X/G�q^�E##�x���c.���hLX!AUv�Z���X��P �h�)�H���?��3F��{Q�%���$�O�j�.oc�|��,o�C*�{�k���9���k�_�w>�a/��{a9������h�y�Y �a �q.X�mkj��#(��>���E���D>�3S�D��;g>5fh�N=�����"�L��l�L�݈�	��dC���e��W�k<��ͣ���t�Qf��w� �Vj�������X�㘝��?��07�O�w�z�osc#F�%�i!#P\�.���/�+��B_p�{��l�a��R]l�z�^C[��ɩ��O7/�c7&��@v�G���qX���{j�\H����q�m
����e�n	��G��/	�,/��kpCӍ��_N��"��]�:xy
`�_[2���(l�����!n������Jg��D�l���@~���)\�Ŭ8�֎�$�v{>�/��x���Xi�Z�lz&R_����>p� ʥ-w�C�Q�,{��	�5��Ҹ1�t���W@:d�i�2�����7�����鵽;
�Ҋ�����%�@p(!Z.��S��6��>pR�ː'�3�V3��?��pe��V���U������?�4�q��C�jouaQ�D	QφӲ&�[���ꉰʾ��l�?L�Z�Z��~�+���"���,h}Yb�wAV������_"������?n�����l�VpL�^���EÏ�1��W4�b�Aft���YR����@f^@� �)�x�4KX�$���L�����tY=��"�{� XkKl:�]|g�ӼP�S\{k��<@>e����.�aB��R���;T܋�Pj͟�k�6<�ͬ�A����z����2�>`^��*b�M;�	�Fuit�'�޽�T��R,��h�%͚�����WQ6�)F^_�YU�����b��'D�;7{I
���1,~5�b����mDdv�)dU������� �;��X��\��3_�c)7&���k������(���<�A�u4��P����2mtQ>El��������Y=g0�b��F�h�:�?�A	L�D���;.:D���i�J���l�����}�1͚5�-U��I��s\_ɵ;>~�7���_�x�������C�+������7X�;�-r.Z��˔�Ј1��8�;EZO~�i�2��G�s\H� ��.����sg���+�E��2�YW#�9Tٌ,B�̚ʔ�x�Ҏ;5���n8D7�!Fp{����q�5y�����o�r�ض�Th���jjy8��ە��uhqk�����ܬ�5�QWҟ�.Ȏ�R+k�8d�!�s��D!�;�K}��B��zM��/BEn���!���w���bp���}��&��z�ߋO��5e�%S�mm�p!�����ۢf��ꧣ^`t࿧�٪5P;�*
wU�2@M�S�6� G�؉���Q£��*��	�ѝHl��Y�~�5��wM�,,2)���f��������.�2![D_	�f.ܲ���0�������jCcS<W�}�n���62�T!�.\(~�EK�4�6`|H����N�ȥ��n?�=��e��3��1����4z�+<�Fݬ\ۛ�;�\�$o�޻P]�o>�bC'��Ae3I�}�Wda��\�i�rF?��g��;��K`WT��!�93�g-��0ѡ���	M�Y,�*2�mZ|�[���V�h�.|9��C���Xoe�����
�\K������dxlz��d�ɩ��a ɺF��K	�r���H������g|��[|.G������7.�)�N�c9���kۙ�+u]�����+GOr�s�I�V$�ku���mo�D�bQ��s�-=��F�4�P3�+�� ���R#EY�Pݩ���9WV��iŮ�߃>Ie��ǡ����h����ھ#0������R	-��8rxM���ɜ���ɚz��E�W��F�'�<)OŐ���Q�\����L�}u�ܬ�di���w��Y3<lAy�����R�����9�@v�7s����5�K�Y�$q��{d�2Xh����P�o=���?��Ӝu3�Ŭ�6ݥ������9��`x:b96�p!��g��g*Q3)TE��U� z N�g}:�u^^8�0���qOe�.p9���Or�����f÷�j��b���<��4�u!��ܸ̇\^�`��jˆjub�"���`��	C3#e�K.{��ڹp���I�80Q�K;���8�S��� N�vcĐ0&��1�ÅӲwFi�ƧWQݬ?GC�Id^�$Tk��V�B��Q*��Z��AFt��^˱��B� g�O-�DFǫK�$��]����@��^%(�i[�Fm��i;�O�RL���Nb4�L��\ɨ��V�u�Og�#�YT����8����7#Z@�!���g�� A�~<�T;�9�-��d9ڥ���r5�.��e"�MDhG��%�N�z�� �Ѕ=*�Uf�%�nC˃4��z$��7u�e���Ϥ�Fr�:
�Ā��H�Z��a��*� ��(=U}��򃣷��,sCh���<|�J-�3�8wr��uܳ�K0ҹ���B���A�]do,j,1e�)0��'��P��95 p�T��p���a^Ĵhmi�G����[����{�'j��Q1ws����4��=Yc��'��)i�UȆmB��Jߪ�Y�+�=K7O�)�&�`��R��ەE䁴1uB)n��t����iQR�{���P�_��*C�,�n��bbҖ�C+5z�o�y$7I8�M�o�i�tw掺\ȅ�xT`ۏ�9;������p%��\6����nZ<�`�wK�S� ��C�1��'1D�ҥ�m�r��Y���b�h�Rj��(�n�b�XV#<�)K)�B��#��u��+���G�x�?~��J�Ew�`���l����K����q���P�WQG��\�7��ﺺ�k=�Sn.�]&t�,oinr}���t�c!	�?g����dd�2kD�>�Y�Pֹ}a�ع1��zǯ�۾�u�"�����K�2�{�9/3������[zt�h90�PD�J�V��ERd���V�A�/��,'c��Õz8�:DJ�����8��Q�g�wtD���+E� �V�����2󿣌���̆wf��N
�a�Zy�s��<������e&+Hgz*f���d����g�O��ϐ�M�����ͫR����P�'�R}Z%ЮS���Lݮ���5��V^wp%*�ty�S���#Q~�9~�fI��-�Pք�g����w��"ب�`.j���ɑ�ǟ>|B��u������o2���F��AM�{�5
,�>��V�=����7H���*|T�Fh)xX$d�Ol5ćSaK�!�� AP	�7���c�i��:�°oJ��b�����9���QV�<���;M�4���_��3R�]���}�Qt�;���+${	�i+�J�h���n���<�P6ߩX�o�v�H��"�����:e�Œh�\��0ly�5���p��/�ϺSV�NUpȜ����7>�4�m���׊�i�f��P��Ț��%��ό��%DDJ��-���;F��Q�,�c-M5i�ǃ;�ei���̒N�0<-1$
�QD#�nm���5µ	�7��@��2BUJ&]`W�ޫ#�Qn����ޔ�I��_�����q�Y2G���ǔ_�DtY�׳������d��X�gC��n���H\.f�n�h?�SH�"�x%4H3��!�'C������A�Hm8�O쾈5������#�2���~� �؞_�$,�A�����9��8HK�����%��'@%��6���;j��N�*Ȕmq#�`�us2q�;�u�fF��"�bv�~���M
�g�UC�l�i�TsK��ֿ>
���zb�������y>��򧒴8Aߏrd$꿻�P��x�2�-�KR���'<����nF�}
�6���c�� ������	gn']|s�}��(ö�[x�������u	Y����.d�����6T�u&f�`���DR��KP���3�1�QM�G�1�r<����gJ��po�Z�zV'�}P&�յMi[(Q�+��$���Fմl�i�����d��QQ}"�3Hd�h���#FCk[�a���*���dQ���xR.�§�l�
�dH�R�Uw�SY��"/8�Y0x ��tl��gqs��Ʌ�<�DO�|57.��y����i����S<҈D�{2���$����y��̞��r�`�	��Ǔ(�4��Z�b��6ݯ�����TZϪ������w�nڇ���:n��C�4ٍ��8{2�Ջ��$bH�b�|ǐ��Eo�X��ԋ>z�L��?�]��#0�4OA����	v����u<y��M2���k��*f��:���9�" �H�s��*�}7�^5���t�eZ�R�B�3���_D���Pv���jH�u.G�+�T3.�i^�;�O�u(BG?-����.��Ԝ�vߞ����Ja�5��H����"��O[�O��9�[np+�.�:��=E�����Т��GX'��;h�B�!sŤ�4�}�h�U��BD#;S��EC�ޡ���9bɰ����r�%�'��~���	h��+`殉%U�v�hhmze�<���܎lƸ��m���S�S�U�Xw�jlv >�/��\l�#�J�gX[l
.S�7x5llW��@X���;䉠�Rԇ���C,�g��6&
�܎���*��ߝ`,�"!�����S��5(��E?�������� L=WM�g>���W3)�ե��$����Y��*��xm�J�1��&��4 �lLzL�tЙ!�o;�A��&"b�z��S� � �J�F��C��C�S!9���~8�~fx��_�@QM�4�#ᓓ�Z�R�lz~;e5�$�
~V+%�;��k��$i�����Z\���~�H�ϒ�[��Yؤ�������Q�j��kbi9��]�3j)�t�j���dϯ7Ooir��EiݧHT�0N5`���V<�8�lB��u��X����Po�,B�n�[�VaX�J�h1����f�w'	��]�M�e��<�pr��g�ƨ(/7(]NZq�/+�2�/�1t�&`����<�:�X�,d�ib��H���$f����R�,6���a�����VF���c���<Vވ�Tӝ���ک�J�O=v����������=a����|j��/�5��y���0b��G0z֪�!���mQE��Ҭ�$_�z(�"���a/t�����Z,� Q��:���}�O�N�+���rw�fio �a��f	�cF��>�9�Sr�
�<���b�t?�i���׸9��Y?\�c��0
9C��9#:��]Lӏ�URGVDdd����4� �x��p�����}��b��Z���Ԫg] ǔ6Lp��[��M���$�5��q�qҖ�)��*�2����蕾حf������o�Xh��{���l��D��݋�c�B1��^��f�����?]�nf0? 9���F9�'(�ōl�S�g?(��W�D�xd��)#��ش�lZř[���h�uJ���h�Š�cO����pP<�\���s�<�����!��)W��Vڟ;����PC�u/W��|�܀�Q�".��x��/�
p�!����g�&��|�	���J�枭��ļ���mTW׊�$�l��=��꼶hc���y��}������|��R��V��4�TgY�+�h���C�Bz��^������!������*�}C$�ݕ��.ns�0r����4�Z�:�6�@7-�VQ;������zC����p� s�Q3�E���HLA�oSM����Ϭ�7�M��u$�5΃B���{{�q�m�%�M��#`���|n6�
Iؔ�:Ŀ�UH����.6�) G�W�i��wm��i���|��W�*�(�{!Aw3�E�/�������6��K'���0Z�@�4[6��Vg����q�ꛛ�O�Ŏ��h
6���݁+�Y'ݽ�e��y�fH��7y�~�*�A��L}ﱓ�n�.���q���*����*�M[�֮K��y����in�%���=�� �`5;�iEqb�p�����p��,�L�v�*
�H�B�VK����m���_^��hݪK�G�x��S0� �f�!�G� u�IcnAV�?��̙�4{�*�X'��ڵ�o�E ��b	T2���t,�m�M���59�\`������P9��fX�k��&ti�`B�0�zE����!#?��(gz}"
�R��(?�ط���8��>Z�ϣ-�at3�YFZL��5�|�Q<D�H�
�s�ѫ����;�w���"l���~��̟Y��v(������A��Xl�hUxզ�>�����|�oe���h��-�Ưu�g��r�u{��2��m��z:�U{��"��3q�㸯�����n@Q*�bؽ��G3vM3��T��@o����x,_{�����z���&���R��n	IG-%�]�>S�(^�s�Y�'��A�&�k�%{�:�E/�1�YW.�-�=��g �.�+�����-,�
e�Г�N)�6�K�6~�-�1���Q�����()�Ԯ���\z�SIX�0+�ԀbCl�o�b�����Nl_fJ�5���bޮ���e�G̔6�iG�v=���<]�A}%?�������W�<y�����ǥb��J�$�!+��a��|I%�J�5��m�B��1�V:gR�2#sU���R)�[�bA�D0�WT�7��tN���>.�����v��@Jc�f,虎n�-��I֡�cuv���89X�"��z�R+�vy��ъ��:���2hyy�����b��s��*�(|<9��;7�M�6��atD��¯�?!�t-��l����[~����pfUk�u�%��s� �\�As�Ȟíu*��f&�}(䩕�$EJ�6q�t�0�ES/)�C
�#Nߖi�������G�e��e�}�P�k�uۈ���B xr����w��/da�/C�2�{�q�V<��k1���\��FG��H��D<��D񪝷�����tbCcP*~�W\��F�!�]_j����7S�cZ9n�X�T�(�T���B�u���GQX#��M��/���A%>٢��/%.o6�F03f�%�her�~�I:�O�w�ay����;q��݁�IX0�	B�4�zt:JLժ=Q� !��`�e�P��ޛ������Yؗv�ւ8�a�l2���QcS�r{X��cǏ����9����Q�Ѿ��T`;Z��N~���w�*;���?\糂��{��6� L�C=�p�߽�iy�ET7��@��*��l8ͷ�ޙ|���|�|[3�H��[t�0��x!������Ϗ(m��%�ܘKHV*=X�H�}],��k@S�<?���R	���iK:`զ1�j�G�M�J��D�P�],��r��A�SC	؍�T�g�a�ty�uU���Ee�Q`_q[�iX���6�������l. ��!.d5�]BG�����^Ժ�,A�N�I;�J���NXp�>G٨vϩjHa&W������Ǳ�c��������3��ucƖ(������"�a�����j�>h�7��j3��ecz;�{��|t�L^�/�>�D���C��9�?_�Ԩ�h�@.��N;��*4_y�J����헕��:>,�Z�.�]a(݁��I��`�;� ��`$[hn�Z�YpBJ�A
�tq���2I�<d߮�m��7}*���F�A��"ci�����n��`D��e0��S��H2�h�{<xi��et�h7�'�����~	����t��#{ �N��g�MØ�z��&��2���.��3 ���S��#�n�|]2,��G��X�hǟ���ڸ�ܖ~3 ���x�N+���%�F1 +w�����F��*f֓���� ����L�ݸi*o������Hf�v&6��7V���2[Z��J�1��3�/��/U�X���2$�g�8���7˘oXM�C��t�K����ǻ�9�V�~���X/O��� ���'�������x}�4�$���N�ja:'	1���Q��y�&��ꖒ�4�c:��P.$>l�P,�f�o��I�ӌM?Y��n��y�7B����g�أ����A�C1oZN����[��W�q�}\C�n�j�����؛Qi�תT�A;,�'Ɋ�\0r�{js���<��K���WL�nk���=����=x+��G�'.K���\��8��(���O�-u��wU�i.{��U+����:4y9}ᗙq��;F������ �<Tc�}ޗ@�
��s�L]���wm�=�ۯ�K���o���@d����^P��n`��k��Py���_��� ���K Ef��C�j��%�a6�t�]��8�}��O8Ձ, M,���~���U�F�%��8A�-�a� ����X��Q��M��X����9�'�Ġ�����U��O�08�t���~�������q�k�3�r�l���g1��#����\(�8�8�������&�6E�}�s|�'��cuC��fv)C��������;��_|t#�JZ�B�P�Ŗ�8s�t��*����%�n�h���u|G�ϣT�bRw�I���h�!��tgg���E�O�.��P�,�0��g��q��Og��V�=b��PiwjD���x���ށ�^����Jb�(xL�hF���T��oÀ���r�7ƨ 4�����?��1jSN���g�d��V�a�ELYY���D�YO*���"B���bv����J\�#g��E$���L'�`���C����1�Z��`���R0�R
�h����:I�]�:���F��"R��Sxu'[>����=�|�����u�|�֖�e�}�7���2�x��j:��	*=3U��yCt���%KG�h�[���+&XH:n��F!e&�A��& �n-��^i(�4NM<MI�-���k�	t�`G.�����BvT�z}A���&�~�EY��Oum��A@E�&�~�Uu%��5��p���ʜ����$/5~���s�0\yg����+�_y�<�Q<l��j��3歌Y�&2c�_� �b[�+=�u��m6ws��s�P\"�4h����Գ���
*�Q��O� �ӡ���f�h����i퀈C�-+�aW����o�D3��I5&�"׌I�wG�*�UZ_�6�@-FN��~M�~hK<�ZߣH�8�up�H}�8G�T�<I�8��L�lC9�|�4#������'32�xͧpg��U��Ҽ��$Ud�Pi��b�)@�=�|�)�hͩ�%���5ԗc7>*��e�@)�[xڞ*�9���Q�� (A��z�B��(�H�R�6~84��b�D0�{���}�@q����+����ͬkO�u����W1�h]���j��=�kXE����1��V�qH���c�q�S+;V�����p�G$�4��������X��������A� k',@�f}3�A���NU`wq����A�D�^�IԾ�뻨kT-KO�M-��F2�8�a�p���pT����;����SI��N�!l��e�;2J>[VFE�O`��@��*l��έA�߷���3g�8@C�9W���X:�ۛ
k���	�MP���)���$kW� �jݑt��(�$Y�����Mטn�P�{�1g�{?_��\^�_D������5�̄i9X3Ž�\��y�@N�ǡ�+�Z���1F$�E�X����6{A��4�� @,����M�����b�P���̲k���<P�����v]g��@2�D�E]}��q'�����y��L��@k��f"�Xۄ$j;��]�_[��s�rX�!����?@ ��v�]>����M��	o�M��V�,���'3w�:�t�#y�A�w��ֽ,�M{di�G��SU��s����\��V,)r�`����ZI�|-K*��i�t�q
�h^�U���G��
���&u}:�P�j����H{�nLv��|�k�3A�i���<f��s]��
�$�q�8.K:��r��$�i�[��;�Y�@���I4�(��,?�N3"��_�X����$�7@`)��ЍH[K�8�' -���C����[��6h��o6�8��s!� ��u_�
<I�=BQX����������7L�ǣ��b�ځex9OL�8���!�^�4U�����ߺ��ͽ`�`݃9��ޔmU���t����7��NPS�8�9���|W���bn�� <��/c'/{K���6�3�	#������`"w�M�Kn11Qk�	�U�J>�n��� o��B�u1H��R�ɒBE�e,�B��}u�����\-��F�P+�Q�W�%�*gt�`��+�7����b�m��9���X��4�ٶ�谉��)������D,,���]&X��JB\�c���j�����^�q`y�igx^�A�%*���%־�wv�S`�������	W�qr��O������8�M�n��/p� �3��Y��K�4�\���Z�w2@�?��)�T��p\�	���ޮ���A��ܫ��X2
MNFI��>��G�o�#�'�ޱ%��������������ӵ3�n
z���j�P0cҴ�h�n��]��Б�B;�=A�}Hl6��T��Z�z���Eӱ��㛯�R@�&�Lo��P�����6��#7s�D0+@�Gb�d��ץ�`�W�n7nd>�=��LH���%^�a:���"����Q�?W3$\87 �"P�)T`�z"i�U��CL���v^�ᛞ)�G��l"���x�T^�좏�[)����۬Mm`�ܬ���5`Zx��d��.P8W�c����vG��&�O�v���?O��*ē�`*�/̫�R��������R�/Z���$��]����)wb|+j��Ԗ#\A�qYs9�G^�5q�Eo��C��'����/ʸ��>�@��31u�ؖ��	�^}���W�3C��H3�&ӓ�F]tf�S�ij�>�?�F�Pg��0�H�O�h�60`]�į4Q�n��9�D��	l��=|�� M�+�&W!����>�*�iYV�a���Ż��l��`6B����7O`diLj�)�sJ�M0���\Fu���%�M��U������'Jګ�6DI(q��pa�2���c�7�� 9�\MV��OU�J����(`lA��MC�f�:�'(�k���VIp��'	���3�U-rI �JN�j��z3]3�o���ְ+#P�jK]c&w�rf����.�Xd* mi6ط?�$���U�=!p�_ԅL� ��`� <��}�q���R�E��H�	Rv��ۼ��m����E�~������a��ਡFVr�!TE�J�������S]�|��t�#�=c9ec�˒�P�w/\e�'7�hXު��cNfr��͛��Li�6��xV�K���}��=]�tsH �M�3���PAq��1���ƍ�Y��QY��:1U����e(c�F�D*W��ֽ�[�
��uU��?��M����]���~�q0�Ĩ��MH�K�,���U�oKa��!�vF]������jܜlAP�mm�ҕ�s<�#���{;��ԉ��"��p�@��i�(����x�AM��+(�m̀�s�is?|��1�x���E��A5?r����a�:wOEc4�v�����t����G?�r���vҏ�s����މy{��)2����IW�!v�t�6�ch�r{\�̛�郚5c?�/<�g���c��\N��ݶ8�VG5�V-Rbɠi�n�×W/�J�yg�����ٓ�Q��z�1��2�i���#'yy���8������a����"�T�D�98R:���}�ʋ�P��]Z?�X�c<K�� o�𵶏VdxR�jziE߲���H{�Y���ԉL�n<�+�P&��e��r<gb���pw�l�[��mL� �$f=$
E2����N�Jx@=�-(�9]h-%S� ��P&-ן��~֮l����b��A��39 �3�i�D(��:�E*'Q�k���#����(k����L��}~���=��;���9����,�����V0⇖��m��j��ad_�۲��:.2λF���'�,e�|�/�tSo�'z'�R�1�v�R�%�n"�13�P{o��]Ay�8[����`��pb�񓫚�\4��i?S��E�O����P�w�b�j�2��S������Er2���j�c ��Α�s%�@����}��C���]�"�r!.C�>�|isv�|�+.�!�ԅ��KE �]��pm���f�6�)k��g2��n��?�J�����Rl`?BL�# ����L���}��8:n�1�˔�D�a@��,�.p
V���n�"�1X)����L�������+L��Y�#�㢭��G�`�0���h�kA������@�/�d��JF��&�˻tcb[#-�{�~D�g�~�IL'%1��h��ҁ��l��5��ݘ��qf.e2R�AX=�;�Yh:U�6�Ϧ19�Q�~�cՒV�TO�,N�� �E�t�K�+D��:���UA#e�	l�qB�$��4�����<2-oe�MOG>�:��(�ʩ~�J���j��צȥsK�A��!�>��-�\ϲ`;<~Cr��i;1�`�c��̃�	~(�)�W35�{7�Uͽ����\G[3�ż~��@85=Ŋ�q���2g����S"I�.�g��!��3�X�������E1<��V��Rn�*�yf�7��ʍŔ]UE%Ymt�tr�(Š
�lB�x�2��}��+��PB� �c�Ě!U!���`��N�
�;+�w�ɓ�'�&!���f7g�8���^{k���J�X:�V�YW�&�wجE~0z\�O� [ �A�yt`������1�7�����O�{��Ҷ���;[��s�e�M���`���¨8x��E?n��%9��k��*�X�����6�ߛ2���WO|�.:��T������Ȧ-&l�����'��>��C��h��'gOS� �*�x�s� ���*��Q��KN�LC1�=�ت_�0������=�=I�%�9k���4�VLÊ��ffgL���^���
�QB�ɽ�rҧ��jTA����V-D�n��,���biN ̇e��j�X$X��@�����<@�ʵ�K�5Zv�siw�R�~��R��b�(=��O�hxZ�چc���&�¢{X��$(������-敱�P\�w%]� ��|L#1�+֗H�Q�Mmė	����-����ʵ�블�3���\���g��o+K��^XQ<�|k�Ӑ�T�Z�������g}�6�����V�ٲ:̼��*�y��g(�������qA�lS��X��b�i^�;��� j�����̸����O=�brk3�s�6~�n���V?� d>�E՛zهd���~�[�q���f�����:c�s�|c�+�z��Q!Tp"��n�*�^��-�X�(�9�&I���rwm�E����׵�j �:�e�H�NM��9��UI^?k���H],
_p���˖��j��P�z�C�
���z=k���1�i��m�h�uf�!�:P��Dd��XS����ۨ`k�ԧM��~9�l�\��'�T'[Ur�rC�!4�, qd���*M�x��!|�8j�?a�w���PC�ɹ��`�w��Q�>8���	�1����PS��^���Oۚ�8�x�cݧ�m�_�iC�$�k	�(��Q���Z��퐻�yx>�=�������*�hW+��y�N���^�1H���=K�X:;�� ��٣�WuGJ�t���.����ك�Mf�l�p}��L� @^�/��EJ�)e�k�u+O��B�H�%y1���U�UpP�ᓓ���D[T?�I{���Ue��G�L��
@�k��l� !m���g���>���$n���[�7�zHW���7�I� ��X��!�F1�q�(c�H���2=�줷����)v�v��1��0\�l�;�<wW�E��A3� ��O�@�[#��V'��dT��Q5����u�9t4|F�E4tÿ��?c�F�v�ɾSH���/�cY�1�lI'�c��4�I�������[��\�%��� ylƓ�Y���gA2�A=�]6W����F�>0#�Yh��Cmh"ô��3�+	��fg�' �&�ۺ��J�k�G���9�
�x��'���'��9A�gؠ%�_䉦��
���qUGS��2�sW���c,p���ɘƩ�9�s�r>F�^�n�J�x���f*g�/��x��T�,��W4�����{5'��1���;x[�c �En���T~i�WU������&� ����=�;#9�u�X��A=�6aOxᛰ`Չ�p<QP������P�FQ�����<V�t�%N�2yT:Lݡ.,(���S�C�F5VhM})� Fǵ=Xy!/��`�{Rd���Am�=����ՠ�)(2}��j��GK��
�s)�^ �;?�Z�7�Ɨf'#{��B���7���s[���3��%��Fl%�#K�'�@mb4(I&���?�F��8'q4+3���;�#f������V�r��)/&�xdZ���=�T8�L�Vq�R�(�{���ߺTi"tM9<�29B�j����(F��ji�XS��fy�!~W'�`z��Ҁ&C=��)��]���#�3 ަg� �4�{eƸ�nBZ�J���&���!�� ���\���W�}&	b.���R�Q/�����:�L��H���I��`�5��K�����[���hL�S��6�#N����0�r�73O����=���"�W]cd��`�Du$���Yk�	EK�	�GQ�^�.�J�ɷ���AM��>��^f�ϰU�ímL:��7�*��v zNhO:��9���a�R�>\��������`D�M$!�Kж~5�-^sk�O�c�H�u�/#S�T�Z�r�6�|ٻvն�͙>�����&�xD6�T6W=�w:�L���ĂI��*��W@I�� ���p�g���_4?~3յbG_ϰ����y�wI�x�8J2z�gc���G���ݟn�\� ~��) ݜ��A����h��O��!Mf�I ���=��~����ʨf�&�����b�g����g���'�R��
�{y��j)t�!Z�-�]n��|���E=l�&�y�j)yfm��N'�����`�l2��v���(4�)(I� ;���p�q��ꄬ�nSJ10���5/��*��|�����g"V�R��s��̧)ｃr��u~���ۀ��74C���t��|��F��iy�[/sʸQ�'���D�t�ي�Vz��-���?[��+�l��1co���wZ�9SD3���V@)��り}~��G�+��	G��d=�z�^�I���+1�����I�)��5zm�#'�C��E�h9Ɂ���K����m�F��џX�(��{@c9{ĕ����ޢ�8q$hgR�!+F��7�B�T��*��eL::;ܗ?uJ{�3���.���AD_��(��v
 �օ�;�yu'"0g(�e=��=a��1�߀��4R7cw��)�A6��N�	;	����V������0�~�b|���IXH�u�N%&��Q��{��V��$0��,|@8#��!Z{����l�M��8�M&+a������b�Xu?�/&�.�T�%s�i�3��;!�>�H�Q�#s'�h6��� s$@Y勄�bh�@�}�[��F� �lWK}PX(ǰ���rl� ��M�%�7�~�~�5z=4G�I�qm`�f7WDw�pF��d�7�S���<�P��/�Qh�Z!�a���xP�jR(A}P qu��(l���2����E����'-X����q^a�WMj�<i�i���$��n%jA�!��f��b�����bW�j�S}�E���M��0w4&�/���r��y��zM~�H��{��t�N:��<�"��˻sFﰒG�/�,�u��"�ĦHě,�aj�u���=i�a�y��O���4hJ�k}Y�v�N{E�6f�2�lt��:͎nX����b� d�C�Aˋ �����9s���ԇj��Z�6�n���1�\Q	c����܄��7�*x(�j9q���3��/������M����F����)�&Lͤ�b���@�������*�Ty-$�^Yˁ<�I�|�7/�'�OP%�t#
��F'SJq���TIZp�:��m����L���/t�DN�|�8���8���k�߳�L����C۱����I���ΧZ	rf�RW4�:iY�f�V�O�o[�z��Ee��c�I�	x1���{���&.%�(��1�W-� �-q�c��$ ����?W�t����&�!P�N�򉎄a�xaS*��j�ݣ�e*ߌ����W�P�F��?��v��<!���hH�Xى��š�j����"{aK�v��4^�l�/M���#��]:��kY�O�.WmΐW å$v������\��6{�J5j��=Gp��Q�0-�ng
�h)R>�6��굿J�)뱊ϫ�s ̪���-�'y�ژs�6α�Izm�,�'��SC<�/��dik����N��l�;�V�B�9CX������H{?aU�H:�2�0�k�pMoԚ\�|<e(Ȥ��pa[��?����I��ol��5]��o��~�%2������!d�|��-3��'BP?��h8>�-D�b�q��b��N��O�W`a�[b"	#�|qGVȭ�f�Y�1=l��f0=�
j�;��5��5��ỷyFw7�^��r�a��¹���*�8p��{�9=�C�NZ��z�d��'9f�sS���>�Q���ڙ-V��?�f�qH�5�痮�~��n�%I_��SEP���b�]/r�M�8sj�$P��l
�@2�!>̰��>9:Q��	U�X�XP���I�c۞�@޵ϧ7�#+
$X¿�m�6Լ��+�c���v�GKh-G8����Q��AZ	�Ief���Xi4���<I�D�^ҙ�[�6X�����,	�=0�����H{����t�2�3��5����։�k��V�[}d��@�5P�B>j���V������C���
������JW@-?X����a�2J�Ke�Μ[���y�����\�������{%���2mP�H�����������-�{G���5��5�ߩ��|��"9W���#�{P���P��e��%t�NAPO����1��u�dS��)ŗ	S�q���c4^J��x ��-����*T�rD����@��m1�׼�L��|b�1�")h��Q-����k'IdA ���l/ӫ��"��y f���ܳ�/�>�J�6p�ڊR�0_��(�{�a=�g��r�;ӥ�sDTx��@�&��#�H^��r�{�!����Jh��t��P����Ų�5������\��ӿN=���ٙ1D�E���s�a��K�}t�q�����عt���w]b@&���l�,�s�9�������& )���\�Qm˂������o�2yM�M����I"�~��LA���d�rvbxEx���i8��)=.2�^���g��3�Ua&�DA���玗�����O;ԅ��˴t5���F�Kb}R1�9�`;t|D�{��'�Km�z,r�1�[BZ5��c�����cg�YK)� hR��:���|�6����v�7i5͏r"c���U�����T�R���j	�yNR�k2Eݫn����fK�Js@��rm�H�>�I��nh���>lw�Lg��Jh�G&�֕�!.Ԓ抳�Q�2o&5�8�(G	N����q��0����8W�h.{�b�Qbu����c[�t��������N#m�a0U���1I �4�7�5=�ۅ^��VP"�l �f i��<���yKX�!�?>j���ўG<����!pE��Y��0�n$��[$��"���K��D�^*�������j��sV����n�Ԩ7MM��SG��_�I�l�LfƇ�Z@�Ǣ��Ti�^��F�;.ఠBp/7�����M����}���t���s�
�������7!�&���gp�f��6;s�
o��׀��ZQy2����tC�3ɭ�߮ n�ϲu�ժd��r�%gp6�ֻ�,�2&I�>)_�3��=�8gjS��T���%kr�b�s,C�E���'�R��`���š.<$�ws��4!Za��j4����y��ྫ���y�Uq%>�����d��C�[�J|Q�f��g��x��P��g�*�],\+4K��L���$��|��.���8+�c͌�h��^8�ޭ�@7���|��xzI�3��~h��z���&��%F���Ʀ��$8;�M))�I�p�E��L�u��P0<��k'A-
rf�O���9���Ԉx�ϕY��2�';�!z<�p�;=�.�� �&C� zHh��V;�zH�ys)+y�������kL����Q�����ԑwX<[T����Ɲ�;�u�~��
����n�MU�ˋ����W~jh�n�y:Ϸ�dYwš����_���\ثեa��b��M�{5R��&��ޭ�̏���)��%�X'^���v><��V�3��f
��z�9X~�����+<�E�N��k�o[���n�JP�;�:w��O�l+!��m]����7�� �1r(�O��@�c���F.>�b��͂Z[}{)¢�����W���W#A�S�����Ueϔ'X�X�����a�/Hn���~� O� t����^PaE/�:ɳ��e�3��w�~y?/�������#�%q�;D�2MJ�4}�HD��tR�~��A.��m����jzsS�}��E���	����9��f��)�'�;��I~"�N�X�*�Jo�
���ӡk��Z�'Ra�|J�'��4�z���N 5�@�G��G���@�F���o���!�yUY��J΀�3w�}��Ra����.�K�ub�^+C�>`Ij��� �J�7 q��H�i7<����إ5'UN9Ɂ[�N��?��6H=G�g��^�~`)�*-�O�	�mVm��>d��B%^˛	��!����<��X�W�~�Z�����oO�jj�s������I[錏+�a<r{�1r�=��S��۴py�x�_�Gb���o_�g�`EɄ���J��U� ���� ��Bᅓ�c���B��T�Q'�P*�}�<��Im���,M��Sv�-�`F�M@�R��˃�,�|6�D�FG������b�ꍉ����#����^8C=G��&��~cCB2%��m^5w�{���ב�ϪfE�Ͱg�BRg�~�n�����@�eݡR��
�׳�h�B�c��1�V���h�r��@*���~�5��P�N}�dHW}���N�l;K6w�5t�rg�pE���-$��w��'W��tc�����'�p���V�����!�ٕ}F�Ċv�?��VC���1����0ѱ̘����>��)�wѭ0+�uaA��ԝ�`�l���U���˞�aimk��S� �廖{7�U�"�P*B
�����9@�@�#ݸcpcnu�b�X������u0*P��s�c�q��3���O���-��h.V�[��j5�}^Bm�:�Z���,��- ���3PP֒Mʎ�5OD4���y�Q`6������]�S�͡�Αo]�5�ӟItq�nD�|`3��a^c����Q��<�D�=���ԷճwÖ��G��z&D'{j;1\xRn�u��<˗����*F�٪wb�������v��tME4?XWOřD�[9#yMT��u74������Ҹ)C��?)��Yޔ�D�?����"�յ�Ɯ���[� ���~eoɮ�b7`��;��N�BخS�k��Q����v �'HF��ZU "�<�_�OH!��{��Ⱥ#a� z$gϡ�L�
�zL�4���7��o�������]�r�E¶�G�Y���k�K��zL���`� ��)�7�P��}b ��
�`�fdQA`_���c�	�D�t�-����eu��� ��>���77��i�	��O ��/,��˷x�:�#2������]˫�����׎�	A�7�c���bC�ۇ�5��6����� �h�q��L�:K
-Ð`(��Hv�w�1_�壏����{}�����54=3h��b�B��䪸�:{U����˫f�k%��E�_� IJj-�1�3��!ζ���T3��eg1�&��3�g��ki>/8�1�њ�#��**�d�+��n0FQBd�A�����	)9�C��)��M1L������ y����ݽ�$~"�f�ח?��DD�fEK0:����Z������{�<��ĝ��� �3�׵d���w
]�:W���wZ���؞�/��hwE�$<XҼ
0'�%�P��; �ħh�%}HWk-���V%�L� �| *ЃyG���`��7օ��0N� �	h{ʓ�jV��Dai�#t��A;jUdz�?�^:��㌛�J�y~ }�.R�!"��������Gȟ�X�2Mlr6�9V�r��vƜ���}H���WKB�N�@�����_�Q}в�;|�)b��M2���_�~E��|/�sK9/x��8���wj�>�'��/?\��*yľA�f�̅�3C1R�m��J{��蕶�Zr��RJY��y�4���G���wy"�z�D6K��'D��[`�2>��+D�ȳ�j]��	���˕��1L;�×�ɘ�1 8���b#��N�KWڸ��av�N��� r���F��b�4��H�� �	8�eR���Ɋn1,,u1b����h������f18�O{�<�R��m���>��H��r>�JhF�y��_���~6}��p�Jiޏ=mA�w�?`�E�������@�3�{Jŵ�`���y�H��-?�-�Q�[u5 ���`Y~;���U}|vSru���pcˌ��-���$��j�'B�\
{�'yl��Ĳ[�98`����������=jB�[&�7(�8e�c2���_ɗ�P5C�2�@�����s�C�3�J;�<x��y
�w����_��&Kq�}��.�6��ڲym��Z�8;4����-�z$-��j�0)Ə��a�����(�\�i��I�U�M]6���Ae�K��H�c���4T��s��8���"3��E�BC��q�#��6�W�n���4�c�$�5ƍqcr�"��pa�%_=�T���K�Jv��f���,*��up��<3ۭ~�r»\�x�G3��O�?/R* ��H]��䪡�y��#ԑ���A4���G�o;��}�f�	��Ʌ�����MF�OT��d1n?D����<Ż��N�m���YU=�^�o����D���H�jĳqM)��g�}���p�~X�S�/���Z�f��u;ؿuƱ</���'��:d��� ä�ˏ����~p|��4#�٧�ҝI����?!O1 X�&7�E�e�(�H�1e\�_�,Y������Ĕ�C]D��ߩ��5�+�jD�`��+wK�e�]w��H"�%w�� K��1n �������^��"�7�LL�8h�I����'`��dǱU�n�|Ĩ`K/��5����A9s�l~R�.˫a�1������;��ǥ4�;Q�)%�C��X[����fr,w� �\��SJ\%��ǖ|l��Ev�=��:����j��ls��ukoH�����^�O"6���t����DX[��Vy ��2��v�;~v��RY��p}ӟA���d3�ׄ���̹7�%��C���WZ�ە�kn�j^�2τ�I\t=��}�M���m�iك}7��⅊��x� C~!{�6m����}J%���9���k�꒗'�����V\��Q��8f�s�oWqA��kfm�����1�r�O���������
C�3�����N�$)D��l����x�4�������,�s���O�-.��&��R����֝�=@B�������X�j��k\hy
�T��N�X%K�u'I[E��"7��t�-bg��3?����T���̯�fr�.;r��zZ����)�����+B�o�:f\�7p�
/�9W�n����Jx &�R}���	�c
Y�j�c���>�G��h=e�+��u�SZ��2H4O��Upc��z�M��-P��I��?�e��>�2�lU��?,��N
��}"�1�'R��y���$�]��t�uXmX�u�LO3z���F��/i3���Ca���U��grq�4�I��x^�}~�q����vn�@=�@�CWT��·����:m�b	)���К$�Q��W4.$��	�h�@�OF tx�zU	���_�[V�i� _��m���~��д$L^i�ȕ-��Uq�d��1�vڰJ�i�i���PP�~m?�cf̏0{��K�(��=ez�t%6�<��=!~�����1t����F�QRv�9cOj|��B@��1�1���t�,.;<��}�e\�Gl��"�K��ma���v�:���FS�\�c_�cW�T����|���<3���o1�����Q�C��..��636��<��H�ϝs�<<��e�Ah�ƞ�,V���%�3�Y\�O�x������-��0���6��X.d)���{�����ߣ�@�ï6�̇��ݵ�{���qb������%]P�M��
�su���vK���=`+p�u���R!_��`���I���_8���B�A?{D�g��/I[��T2!K����"�s%(o�� �����d�ud��.�}�3��'.� �F����8<��7���v;G~����i���B�ihs�h� ��z�	��Ly�W/,�4B@�0p 'W��� (t}b5"��1���yGW���{/�?�#��g�)8lM���>��	�ﵸ�K�X�a����I�lZG��c4�hv�5�<�O�:��wm6�W�_�.�z]���[浧�F>� %��!F�Dʹ���-d<�TK�l٤�-"ޓ���F��47����$y�<%n�i����ZV�\mY�ip%�S).v��<n4X�ꥵ��ӣ�7 ���[�~��#�73[Ie���C�Pr��f��C$;Ck�������4hh����{�B@�Y�����pSj�6�_gJ敝m�ɚi���O�r��#.	�z:K0
�v�	�D��':�JB֎J
y��̄B��E�[ND��왗���¬9�����C�zwd���Ytd"�����������N��$��&i�{qh�¤��TA~7Rf��2ƷdS���AQ�[���!lI�vƤ:U�{��/�����<I�>y׹�%�����3\#`���kG���v��>S�K��+��9Kyi��0��m�X^��J����ֶI��%�e��_.�2#(�i	���Vd/�k�|��M����[r���� N�j)Q��*�'�]#�q.���6Z����-ij����F/A�ڰ�{3���%����f�!����H<�^ّZ��Rp�Z���Hf�DX�3���\>z?ﻄ���X+��a�IW�a����%a
.����X�*`R&����ׂqwW���w^��ߴ� ��3��B*&��@	J.g�zi(7e%2��3��ɳ�1���B�ء~*�L�}T���IfK� �|����QnéY�W�t*�]O����Ё��A�<A�����J׫�g�x&�1�U�-c���>(ƺ���6�Ӻ2CЪ���=X�O��tͯFA�:' �~�.�O�	*�E�u]�Nl.NP�9���L��O�9ң�P�@�E�N�S���#��^W��&Ki�W2Z��2��y�f`y�LQ Hr��XÇ���nz'H�M��WlRO�ƕ��u�'K�ѱ߳�
���9��f������m�����C�G�/��\��|դ�v���uBaTSV��G����2k�Լ�H�`f�-��D֎�`�K��3~BC��D�%�$em`�2B��f'�4
�uJڻ�( 9&�#�h*c*r�
'e��'�����]��$�A7iFd�yf-S)�πpNU3�r�5>�!\H��a�cwI�Lf�$ ��#0[��<��Ѐ�qP!A�t�Ng����=���;-C���.#>�g��'G��$�%��;��'�X%ڽ:�>^o\ �vΨ:RUl��h �7�J��1�r�O��D"Y�^�٥Jp�F����Z��,pKn�?���p6\���-�?,'�����c��,fƿ;Y1ay� /��|(2rR�q����^u]Ҭȷ��M'bx�3ŏ�r�Dƒ���\:�ܬ�f��g9�#�������f��dZ��'�U��ܤm�K��`�@�i������p�1o�s�h��u�����&z�S��+� ,j�Na�Ԇ���LM����և~��E{?7�~
���?l����j��{��о%�{��_�����/�k������U����ml�]��+��ԥ���y�/�wv��Y��m�(��3����Q��~�xKUv\��2w����]���s�r��瀠���ޕ�x�g�-����<?��u���^�E�lN2
a��ֽO�|%��T���%�+��\[)K`p�#�jrD��`]���Pj��q����#\� �����}���^�~��w�����y��]�(ɺw0��,/g�b���<�{TM��p�'�eu'�7��[H6��z��H��V	`?d�����F⽂Ni��xMf�)�C����,�G&Yο�"<n,ov]U^]�s��"
T'f�*h,�Ve%��������.O�RW����I����wN��=��F��k���ؑ��*�h[�n<Ӻ��%\"���4&�������
+�uO���!u��
�	�3�D�3���:jM���V�{?�w��z�;�5��O �A�Wވ�2�(����rQ��̡�x�D�Ⱦ�R=���� �����m�nȁ���tp�(��/b���X���X�H���u) m���bDmd��ꫬELŦ��ӹ� (+�1���y4���G;��/��eR䱓n�D	��L�e��XB�
⏉+��������/t��* �A�zZ*[���<E�W�A]�g;�O�X����ʇ�q�GN���#lulX�S�$7RǗ��ya��E����,Ê��X�%%E�Ǜա,�� ~,���w��4rj$7��v�M�g�~S2ǚ�,#�t��s�f\Z}4+�@�Ĥm��z���<�������7؈"/������
�7���l��������j���	�Jw0��-D�M���p�����6:5�9w�
wv$eT�ᝣ�R"���Z�{@�L�P��kypY.��O�g�B�1=���w�`Y��Hb��N4X���{��e��V��c��+���zk0[��R�����M#��FBy�߫�+=i����O%��s�v����s	�Aqlo1�	�D0�f��0}���gqb�ՐRTW.��'�23�����F�\R2Վ��̿��̥��z�~�`��ƴ�ĕ! �d�	�L>B���/A;\����(]U��C5�Z�i�đ��zL
��ۖk�E�?��:��W�`�7H�~|R�=H���A��1!�6�!	���@�\Yec�����2��>%@��g�$n[#2�@+��wGfS�?!:���6π�¸�#76��"
��xq�'�v����E�����-�ҏ��
�{���-�j�9k}#`�o���}fE�u^�t��Ho�׃��h��3v�K�u�`������T	S���E=�a�ޔr���4�����T	F��R\E�Q�_�Q.4� k_h/�	 {�I��>=@����h�!��7�P��Fk�Q�^f�Z���pWe��y/M�K2��7��Q� D����p�Ԭ�# �ċn��Ӈ䴒���߁��À��r���@���J�"ށ���d��J�`j����S,������'�n��B_Y�L%��%o�u2���%,�X.�y���Bc`�OYk�L����T��M�y۲"C�hإUH�_����S>E%�NǠ#�F�
f�ܚ�n������ERC�뙊g<��PI�� ��}�� �rV�7��3X�x�T����_��ө�LM��Ԗ��9Q� �ر�������7�ƀx�� �Uڣ����MO���&b�<{J_ԠJ%�M{ �:�P(Bp�P%lQ5\�ͫ4���TՏ�/v�#?��P82=hm=�7. �>Hp/��K�YECɈ�[4��4>ڣB�4,�[$�d�u�=�������P�k젂n��C	��o������g9m����r+#8G�gnYz�!]ib�?��Q%[�01����֨����-�wS�
�PY��箬d���+a(�|��Hu)�\�B��ϸ�mA� ,>̎<zv;�ؚY �k�W�3�������r�#���͏���T������
�/@y�F/��8q����=wMO��n�	l�ʄ����R��2Nu찝�L�I�dPp��Y�]�C���=!ݺ�ǔ�,rX��������9�j`%�7]��+4T!j�m^��Ь��:)K����N�d���i\�ߏtMc�1���V��>�-[$�<b�N�=x�iWI�Q�$>t4��!�v�xm<���	ܸ�C�7| 1�M`���(�g�؛Q^��	R-�4��f=�0���ʒ���(u�*����Pf�V��C����ƃ�y�����W��L\���2tNw��ӏ�b�Q�|B�N��GC�!�n��:^e׈���x�}'�{�,gR�j��+�����f�6�aB̰@o���p?%YY��p4z�#�PMnI�R#j �;V�w�����K&�n�sb�٧��_�XXpjq�0����Ac'��X�kɩ�f�g�)�cqܒ䁃�}Ȫ&*h}�����b=���]���b鱉`�]v6�PJ�;U�d"?(��5CC��|��KQ�^j.J5��|/_�|ZHpq��3����N�Vt���D�������֬<��Ą涪�(7�==��ȕ�+��܀:'M�Z5�-�K�Am�.U_�,�%��	0J����3;N�(�3^�*��W��!��{�L����y)���=AL���e���Y��2��k.A�)�3[OE�,�d����w�K{w5������N,z����I�mײv|��z	����(��Y_L��)�e�J3Z��T�SU\�����;�uݭ{�Yȝ{.���c\Y�� x�6�iE�
M�Ip���tK�gM+Pz7��i���q��W��i�t/�XqƲ2��z}k_N0��`�`�z_�ԭ�L"�8�}�:���:}�I �y-�-��Ti����h�d����@�� ����B&ـ����JZ��zgNM���A�F����t�7I�Q:<�n�9T�ɜ-����-J���g�����{'S����^2w����>X����ƀ�`�d*�F��q=-嶶?��58�=�!���4�(9�y�N���Q�V��?+��Y�T�
�ʐOw���8� R�{�/�HM?�tN�x�`��y�@�0	}Ǵ/s�����X�����9�_�>X(����H��#�iG���W Z�k1��7�F�{���wa��8- 8r?<�h��Q�Aʽ6h��L�/�&�������)� }4ٯ�������D�l��1�!�9��T#��T�dN��2�*���b��Q��_�ׄ%�U�G�Xq��Ɓ�k���vW�ظ����)-����7������hmsO#F���@����g�D!�=F9���(�F'�[�1U�ě���I�8�{Ν/���$)�t���g���� K�� �'�g:]�K���<�F�1E�����{�)hy� 8�.��� ����x��!�'Gk�B�s@�,��QvTq]�i�*�:8�$@��WAK�  ��1ۘ������g��.L���D]e~%���6��O��E���iX�݅�O1�`�39����Rx	�H�HO�%q#���W�[����A`L"�k���IEk���+=�g9`� <�1�h�:f"��0�EA9�P#3 G�U��B�d;��&y&X^�wj.A�{��g1����`ـT.ufH�$����sǅ	-E���\S�ַ�Ar�O������k̵^���h�B *�֑������XjJ$�e�J#����Z1[
��lWI�͖2��<]W�ۭ��!�wI�����Dn�K�06�P��8H�g�n��0�/��t�mn�Y<�G�@�0G�Y8oH��-�Qw�fb;�u�J[N�W�ihwi���!�VЙ�}3A9��W�u�+s��e�a�r��*5�F����?�r�<7Tj������w��f>{3ʤ�cL��Xmn]CA_�
�� =�zz&hm��2}���ã�+9���m��T��w���%�����?�����KA`��ǝ��;m�|�ʛ�$�*S��#up���i{I_�.~��M�kD�t�E5W����D@) Gu?$Q�zשI7	,L��e��1��������yFnZ>��[!0��u�;a�ӯ.-���Ĥ���F�+��ͼj[�XG� ��Z����K�����w��)U�`��IM�#�io���n���5B�HۈEhp����I`B&_��\�a��]���B�|^�"�H8���X�n/@�\#�� Z��N�xܼ�b�� �����C5ep?n�2Ԧ�j^o����	���g��*2x��=fj�\0nE��h*��p�y��5204{�p΀[0?X��f��#	�]}k��A>�����z5�䳠��G,탡)�W�:�[���5D�_���գf��psW����L�3�3�-��xu�>� \)�U����5$0����9`֐.�*�UG���ep�`"��f�q�l��s�����F�e��M��[-�ٶ�<��:�.[G����ra����RpRk*(��;m�>nPE���:�+F0��<�_<c{w	�A�F�M�"<������/�C�R�Q����ڣ�K �֠�?�%u�5��E<T��T��%�B�f	׾V�1\�L��'���ˡ$�W��+aE�䥣V�9N�eN���"ˡwhxה	�O0l�?��!jR��oɌ�I.����)_�xq^��X�0�)H1[6J�4�O����`��#���ho=1�Q�;����R��S0�
�� D�?�C&�x��N���r&A2+SG�3�&�i�,d���H���"�7k\8
{hU^��<c1�+��j�`�Pɠ��˶_{�K�N�)�@� ��6��Q�{�@�ӡ�'֖LQ x��Y��sk��Г�`����y�[r�qP��O
hRO�"�^��F]��p�#-u�Fo���P�ږ&>���V�(t��l%��uy��&f!�rc�yL�G4����~��la/��yc��9��$fW,^֤_W����N���Z����Yiy�j�q�����v��ǦK�D	\c.'��], �ts$��R�Ѭ�;�U�j��O��њ�@#U�ۋ4���|�^"]4�S-~��YW�"�&.v��[O�2���=�2�M/c�y�n�W]�[������kÁ����.���$Ԛy�&�Wq��f?�����l�!gM�aH��6��h粢D�Œ��)Y=����q�Ho��i��q�E� dO`��3͒\Fe1���n�yA�s}�^��Ĕ� �-�V���f�`�Eޢ�h�qj�Z�.H����)f�X��I$y�T�<�.z2A�*
��݈�}\��J�W������2�H��4a��U��_�j&;�b4�7;ar�f�r��Bsd�Ip����^"�~���[xbXd�L�z߿�i�(��z��f��21r���Wɳ�TկC_.*�+�'���u
c�۴�O"5t�>���D�Q�؋v���֧��\a�)�u��,����05�Z�=�������Rïk�T��\X�ʗ��w$���xO�3�J�F��X`�`�j�ֲ)�O�ۥ)��R�q��r&������:]MJя_�O�G\�k#K����L�"�P�����iy�N�Q?'	e�Z<:��<hD�H�M�D'�@������((��\�.�Pb�}��AqƏx�B�L�R$p�q&|n��}U1%�A0�,q��tQ�����U"p��HA�H��������q��k�и��F���\��S6Ҷ(ZeHl�)�^p��j�f�*��}t]�?��Aϊ���qѲ��_K����=w���R�j]j�� ``�0���=1ӳ[C��+Y���
�ﹱ�V�7�f���u������sz���L��D���.x.c�yY*���{7��vW<�����X!�@k	E('X�?�h�մ��H2�I��f6Q��u��ʘ2C7��S�M��>��iߟC��V做_�R���
����b��R�<��wun��R8%~U�aD��J[/ף�賁楲��1�R�@��Ȟ��<<����ݒV�Y�@�M�����Gg\�{o���9\��'�A�3�\�5�ܰA�jA�Kź)3?�x��굍�]�_x�'�v[�KĲtsz�N��vU�����ϋ�Ճ�[b��0A�w��T��
Sz
���] ���$��"��,�~���m��vou�[�ڙY>�Au�����~A�n	0#�Y����`i���	Y|�V�
yZ�`s�����7懛%ω:�
k^!A2�{c"TJ����zw�Dq�|°�րX�����6�"ځ3�Y��d��)r��!1��#��N�ߢ=�X�~�~�4�J�R����ֻ���q�WM�w�,R�����	�����T �<I�rA��s<��!��s�a|Gv���yap�u/���8qy���+a�?.�2�9��R�v�� ��O���;��M�!�.^G�j�V	�����O2����ŕ�|'{��ȇ��y"�jI�aM,�ؽ�~R��=k��Q;���x���~��;(�cl6>�W�F0�6��R��ɇ�p�+��`%\�@��mk1Ⱦ!+��u��k��P���favlo�i��$�6��P�f�Y�a�G��B�m�T�㠒�
'��8.^Ck����Ce�ҡ4RK��7eyu�s���Q����J�C�mH�/���5Q�>쒰���E2_�͔�X0��.�� �Y(j�҉�	33�O�v.�]�W�0Ўa3{f�������q�(�d�ڊqo�-`蕣U��vaM��>E�4��� �{��.�K��lb�0X�f�,E�8�����P7�����TZ�(E�P���ޫ����R�Oa�]��:�o�k�aLa��b��ܼO�5uC<@Ч��x�*3��*��>9�`$��=.�I�n�-"����<!���5p�7���*��Z�0�N����Z��[y����D@�!l��r�"���q��A�N��]zՀZ	�t��Z; �(�'9%��%X������"G,"M־�P����k|1�:$��5���o��K�^��Ϧ|�h˅v �Kn�LTH�^�
/T�we,+3y+�v)"wW����@,X,M�Zg@ޏ�?����Ze�w�m�����D�YI�������f���m�����M ��#�$NA@����sNg�ő _|V	�Z��a��1��A�#�4�	�<>-�
!�4�:�d.ۿ���q���Ѝ��B��.��SpB8�t�s���kYC��C[yb���/p��=5����%����8�z�9-�9�$�:����>-���{��qp�-0/s�@T+�!���X�+�����gr
�\�%pFW�����!�]�����X�����Wϴsh�<�\��f6�mt3p|8��g��8d�	gRT�邝�e����!�	2�Ԧ��ծ�����ى�Ec]2�w]Cc�n��#����|^_�x��3�����E�%@� SƁ�R�*�{[.zد�ڧ�=5\)�r�S,vU�8�ۊ��VI�6�^�e��c��L~���*��P.kg6y����^���T/ຶ>p'O�X��3���9�c6���v�����&�!��0�V���| 4L[���lȪ��C��t|��Z��}vmKB���������4�S�����O��H5�Z�.����]�,_/N�v!(������_I�����4�4G�Q�6��'g�HIwr�t�Z^����s�MIFʅof��tWT�h�%/4嚞cZ|BY/�w`�^ܹ$`�W�h���􏾤�H�y%R���'����r�H�V`O�dF|��q���� �a�J�{q���y�5 =�����{$��eV7v=�tk"�[\�4���
�,�(��NO���'�Ѳ6`����h=]��ڷ�5����]�;��wě�//�q���f�M����Z��m��Zm7q5����kN�T@oC�],S������,��t�4���gla�`�a���Wⵋ����]�Pr�u?���M�9�C��6܂Z�=h�I-�"$U���(߅@:`���o���V�_l0���|��E�lǭ�'x)��ݧS	�^��K��yKΘ+	���Q����'����Ƣ��G죱�����%�����I8��5�J.����޹KW���ڡ~�yǘ�_!	܃.�ɉZn�^��D�)�A�Z�=,�n��>�$mqR��N�:����l�rP��E5 \��t�����1ۊb�\~~U��,⢉Kw��ǩ��S�cg~��?�Ӂ�g����ﴄ�x�\Pk����7�{o	 ��]?��m��tö����%ǿcp&+��qWe���	E;r���D�*R_��U�6�b�!�{e'_��T Up�2YL3���t�g�J%l%ݛ���"�R%�!�����І�O&��ͳ���& \��u������@�F�0\�,1ʏ[��ls���@dZL�T�$_W�SiS]:])�c��/���|�9��FK��3;�mrO������\D0ǪF� ��B��
�2I��#�`��^U�+:���s�	��~�k���邎m]����9R�P-�QKTLڦ���Sl�B�o�(���\kT�`���Ҭ�Bp�n�`��O������T�`�]��o�YɎ%w������Hk�i����"0�j��<U	"G�2��A��a'4 �B�����4�w���D�o�<L#�?[C�0���'��#��}�gv�E�T�B�/@�!���Œ6����;�Dz�Pji��c�1��=�F,��0�M�_�(rb��"��!=����1�"�x���^�f�fT���H����wL��k�B���78��G�8:8o&��=�ؘ�I����bj�b?�b�� �9��,~l��l��&����L�l�o�qӑ���yi�Z�`�ŬCp���:~�ۤkKs����E11��&�U2���]����b��^�Q�%AnwѮ짱����~	�h8G�t���O!M���,p��&p�`�Q���!Y�؝Yk���-G�kA�j�����Sv�W�8��kL��Gb&N���Y���wP� _!��E��Sl���	HYv�H�j��W�	��m�6�r�B�%ٷ�v}�4թC����~�ǌ��p.����p�(��_�\�Ѩ��'��ŗĵ�4=���Iܟ���[�Q��OWL�W�ڿt��Yx9	C>���;�� Pm��uq*�?t�Ggrs��D3�dfB���Yd����×R��ʺa^�̄}�c�7"!-R�3�b뒰u���:5P����<o����Z����P$r�Y'�{�Sq��0/�@���'�S/5,LA�?�f�B�+j*=]h�;e�>P���>\�b��m���ؘ
�����@�U7gF���qٮ��ZI��c��Ĺ�zP&�/��M�PU�fs�����g�{t�Q ����\��Bz��eѠZy$kT!D5FQ�p�xV[���,��d)�_JK��`I3";k�����j%�������=����i;�)�U>�Iw=��p�O)�
�`�TI���1�+� ��$+09��Q�����Ƞ��ԥ������1�Eu;��R{(�,K��-��,����F�����"MZ�"��[�u��I�6���t�<�6L�^+��d=h^�_��DH�~W�GS����S�܂�U�1o�I��vȢ$D9+���$�{�h�(�uƪ�j����V�-�<i0|D�9�H�ř��ڜ�Wh��G����|����ί��Fb�T�/ʒ��qZg��� <YFrf9��2U��~j�$��l��0�.N� /��VNR��Q��c�T\�����e�3�
r�i��dV��B����76��h�{�h>L|*M�8�b�xK/�n�̽���Tܮ��&LK�z�@��jn�7(ZF���MQxoK�)�WG ��o�>Ǵ ��G���'�2�"z����\����[M��r��g����y�\�w)� i� &1;��y?	8JF���KQr^����T��Y�՛i_�&}���S�qŁ�gK��h�k1+y��T��pO�ǂ�l���E0�N���pK� �����ðз��}6]���2�BPj`��Mk�v�f���e� �Cר�a��x/Ԣ{Ȣ^����H	$Ω9K��0���>���Vo�H�`T�ch�,��CIx�F�U�X��k������7�5�<r{it擐���R5�{�q֓yN�QI��94��ymSC(�qWs>3�Y��Cm�!��.��ee�gU�t�;�lɡ�u��m���z��H��vo�
[lq��c3Ya�����.���FO��-�t�Q�֒vL��{�")����G�Y�\�`?��;��xfs�^^q�Y�k�*���V���bZ����.f5\�R:'�v_w�p�Fb��&8��v �u��`Ak� �����x,�w=���4p��Y
��q��*�"x�Z_w���Ї���KG����F[�ߗ�	���j �u�5�QdN��.l�?P��)��Q!R6-�>A����O	T�s�<�}U��3����6�|�
��12s�&+����ٸsl��GI�[<>���8��r�Jǟ)��,��;_]N�VO�;�,��� Y�:�o5�1�*��,F�4z̛�bz����aٜ������H:שrsEzK-��i�yc�`qJ�E�/_�h��G*�?CB�l�K|�sgW�>���(��y@�iOp0Ȭ�&�[��G�D������b8Yy�n�S�M�/I�,�)���<S[[�eDO�E���Y%�xf �oP�&�L�c���QQn�r"!�WKPmA�f-Hyܮ��C����AN^-ZC�\.������o�O��|���k��i�.R�4�:}�AK�%�Xe����	a��K�t��鍩B��`��n�'��X����[:���E�S����f\�o�>����q�^�f"�ӌ�3�E�ib�mP�K�=5�Ů�uT��3姳�v�j�PCz���g�詃��/�hՑ���1m��2�/�G[����dwJ��VV1��H�N�@}eΩ����V�cV�O����=���-��#9\��LZ�'3�~��N'�i{��68n�Qd�*l��䄥�"�u��6z�� $x	�ڬ�~5�T��kr�T�a߅Q�w��_ϩ�p5��u�}�%]�#K��ƅ1a��mȖ��?L�f����C9�{�[7�������I�OS ��B�MU�H#���=�t+���v����=f&O{�]J_FG�)��!O� ���`ڇ�@ ��{�T�T`��`:V��о �@�����m�s���Ӂm�r3�|�}'�f�����c$��)�3Ul7STȗ��HǴ^1�a>��`�� �i̇������-f�+y���Y�Q?J���o�������TL�
�RG?�֚�D=9\V��f��*l���],}&-ο�d^�@+�1`{t�
�_�si��������б��?4�h���N��^��(�p�K�2�p&H��XP��&X�x�h�'|��pl�#�\VĦM��c�_{'ǣ8����2��b!N
��yvYnIA@#�OငݰT�K~{ ��ڱ��=�Ռ?g��8�7h���N�GL;P�JF�V?�W���v_�l�.>b�'��za�JR�(�߂&w:�#�V�.6 ���]W���_�9l_5��=��m	T��U�\�_sJ����2��ܶ׃�zT�M���)n���%l�ߩe!0�����r�_��R�M5*�u	���v���d��6���!9�f�GEୈŎ� ���C�Q��%פ�ꎅ8�]��eT2"�DHn_+t�a�A�̫���pr��ɤ�Z#��n�<E��5'ɉw���(�`����2u�7o��.b���iy�<"!���v��"b��Yh����v�@n�Z����f��]�����?"����	qr�-̍��d�~h�Һ_���M^�-3�Uӈv7)�|�qwW�9~{ƳL��._�=���9�q�$���"&�e;=�Pw��~Tk�(,�X�d||�2Z+�>��*�aNjM�y��r2
�/<�$�e|$��ہG$u7W^�^���P�n�#7s0���1�u!�{@cv[p&̌d[�x6O�Э�� ��v��s�P����\:�'��O-���y���<&:օ�����A��ɘ�kD�1�c�M��k �O�.��Ԕ���+~� '�t���bN���ۃ�MwCJ��>le�?�8z�����5`3�l�H�N�&��]�
���Z�`�`���Qb�6o%�A�B���KR�x� Iڦnъ�X�a�nA�����#�e8�|,�����mJ_܇ͮ7�J��T�@���H��RO�:����.oU<��\Cع*��K��KX-S*��@w�P��V;���x;(����Z7h���!�`��t7PI0ų45H���nK�o��\R+�*�Z�~��{�Xn��]�L�%�U˷���&�IC%�����+=^צVj��F���QGviz�>//������ۋA�?3=���^��(��-�ʩ�_�p;�݉�~�Y���W�'5ĢZ�N@3�F>5+A�y��?��P�̙[��S����KU���`
���-:ǝr�_����lo�bpn�!
B��I2��S�k]�O��ם���z+��1?��\�`d\�E����Y�M������;��x������_H9����i~���5�9t9��� Q�R>�-�����|�l�����e��h%�:������4��c{�Չ�t+�t�;�Щ9�����T}?��r�جz�/�joq�������O��P�t-ț�����"u[��ݲ�� ����1��lDE��TZ��)6�x�b�<]�룅��ɺ�O|�~ WB�{;ĝ����SW�a���Y���V�����mP�k%>'J	y�Tq�yCK��`�xpv���;x��w\B���׷ɁB�(�A�����@wv�,7V�#uX��	+-A��R�v|�eo�RKO��c�w�����`˚G�g4CؒC�����L��%j@3$^,g���+����3U{���_����Cy����"U�h���^�(���/��VÂ;6+��j�$b��?�	-�ۗ���hp���j�n%�]������^�i��5�@�'�<X<�w+ڹ��w�Ap�2���I�Y�F�KfI�n��Ɋ�~,f>����'�wH�Y9��l\i���#��~2��)̚�G�!7��`�CDXji;a��#� �^�uF�6�\ws����&W���ivV��\撫t�,��<���=�
y���cO�>� _�K��%�#u�@���$M���3�����u���Y�C3���_��Di�������b%9f����NGE������$E�ɱ('T1/N8Uל-?i�t˯mk�jB�$��)���m��$��m�e��7j8rgE9kt[�Į�H���D]���hh[������ә��̥d�{/`%z�#bل�_���}��0��Kn�'~�^ОNʝ'��$���w�R�J�SF�uo��#l�R���x�J]3�=z�p�Nx���8�1mm�x����h�#�'�p��S(���4�����Ե�ԟ��p�+ޖȥS�
��w�s���4<a�uJ�S)c���hG��R(�hgl��]����g/��g�zA[{��X�\�P�5�%�$�l�h�=2��F����!A�rŕ|�Y��0:-��*^�	��Ơ*�q=~B�k�΅�����Έ���`��~7u'�9�z�bz�Fm����+i������k;�3s�Y!�yU�!E��z$Կ��,6��p��ک~ �

ۈVX)�z���w���%��A{U띲��M�>$�x]|�<�{��:׊�i<���@�pڄh�m�VY�t�%=.��R�a9T��@��B@��Gt瓘d��NS�Bɮ̈��{4�{6�Ň;_��)�.��
~�b�(����8'�8 q��뼊�E�R�T������&�»�>S`�E��hI@�^7R�h�L��ob�s��f�Kv�	�S��!�xn�[�gYT���A�����B�C�D�1R1��9�Ͱ�6� �T��q�_��7��T-c�G�T��bnWHZ���h+}��6����q��p�-S��Y(	e��KZ��̻8J�˩8�I� V�q+�$�Gw��d�i�e�}9�Ċ�v�����+�~Z2S
������n��m�'��?�,�
0���g�3ޖ�x~��G�i;��w���ք����pE僥M���rK2�:L�(�~@���
��}�mT��|`ǣ�K�8�VAR����Su1�Ø	�1�P�:��qK����<}A�[i�4C#-U�_�7՟�Cڡ}�ě���
'OJ|&���hFˑO��*���!K�����:>)v��z��PD%V>	�s/�p
�ʪf/t��j5&����ް�i��wY�<laY�o����ĄXb3 �2S�F�T�����s�x@�=2YCڐ��	Fg�@���7y
���w:H�!h�}����r��Y���@P7��2�N�6tb��*�*^���OH��f�R����^�ox�v'��m����'����+m��\�w�u�p^�I���ĉ�=���������	�)�}��b_kI4��5ȯ�"�P�V'��V�P�0��d,]��0S*��DC�������s?��@<��Hv`F�A��hB��O��K[q�Wδ=�����=S�,���^�� 3���>�rDͽI��`��GjAOf���#������3 y���΋_���!���A��W:��V׽�/4�DE����q./=��3�ƪBz��C#rB5���B�vM@	AІ���$�3�Q<`����:�\|n���M-��dö��s��y�w�;���5u�����Y.��뺮QQ����JPJ2RC��0yt5�Sn�39yp���|3�C�䝹O���.ޞ"�Sc�KT���{�ף-�].�����"��G?dKr��\��S
~�lh0�)�v8�e�\G������	�2���Ҽ�]G��,�_R'�#|9#�BNƳ$�^1�ɲ��f0�lFV@�=-�ϾX)}�7�Y!�d����+d�SÚ�R��.�*W ��K���j��ہ�w�	0�/Bc����ݺH#��o�P�o��1LtΓ2�\�x����A�@GN�л����m�z���A�_v4q=ӗ�a�0�Y{H�F�w���{��҇(��.q��cR.FS�NO�i�d�,�<o���U9��p��#�rY�NzOj"��U�brՍd�����6���~�+Xq29��!�)N�7���g�,��&�¿��ǚ3��S�	�	���͂3d�S�)�b@e�v-Z�_�&H�
�}�U���dW���d3��ٗ���,X)W��=	uG�oC���S���3Z%���N�l�E� ����~q;xr_.'�����P,)����q^Z�~,0ۼ�}��gC~%���@������%A,��{�`N��<�ĭ���!n䀉���(.C���ܬ2܀Yd�f7^��'��z���:�yr�` ���9�I�0kN���������V�[����Ҏ�[p@1�7�G=��1��g��_9���!<����Ђ�����5y~F�u�:﹊�g�8��X��J
iR1&zm�l�h+6
�lf,�<��ԙS�1��+Tn2狫��ϭu�f͞�u�߈7=q�T�9�]�#� �Er�Fh, �$��l28F��ll�ߕ�����=uن\�rH?�qsP��~{߬F�1^ɻr.���r�N�$X9��@������e����ʆ*�7���n4�*+A�六����˰��K��2��p�5~ի�S~��ϲ�5���}��A�s9Pj� �@O���7�4�>:mfy���O� $̎�8;��I&��'��ӟ�c�v�ox/<�(���V�"ovu �/6@�s�~��ə*��� it�V��#rQ��1��a�{S?"�v����0L�y���V�֒���oI�a+�އ�܅rH�����W^~�N�|�	���P�&F<F&��[Չ�f�N���F��*�1��=� �`�Zef�����7xX%nt>f��=�OjBoT+/]N��«��ehSK-�H�uH�~��$=�e�eG1b�̪�[�,��`� ��7�)�P�{?a
�O���1D/�w��K)Zٙ��w�_�2g|	!���<�	�M��׆������>��B�L��`���n� p���[�v�PXZIF���}������r)䁏E�
����9�� Ԓ����*���7ƱDQ}�S�{��/Y
������b�.��D�n�>Je����k�W��Ku��c}�3}���h��g��n��I�ӧy,��XJ#�����$�f�g?ޝ���
eD��61�����e߹Ӌ���s�Bȟ���#h�(u���O��9�GT�#T�U�'��ºV)/ D-��O�J�ƫrަ<��P���Xw.�S��h����QA�`3��l��Aံ��$�P��
����o��E��4E*�o����!�����O(��1?��J[�I-#w�����3ֲ�3E���ٟ�8�W���A�,1:��N̹vƣ� ��]믊3����˭�������Q}M��혝Q)A�?&�N'��4ޥ�x��ȥ�=׊R}�D��y(�tZ��þ���5����v@�#�*t���~�Ք�l�
����kF�P�o�� ��֨�V�l������&�f<���I ���]�D���W�-fH��[zum��T�B[q��������V�)�H#� �l��4.���q
��+�#�h(M%��a��X`�a���P1~�L��(`j%P����á�|�(N����T۴�2�g2+v6�<�L�eGH�O�����(Α*�2{2����ώ(�!��M�����X���{cLV�ތ3��̆��]��>�:�Rdh_�ˬ�tB�-����?��P�lw���ȬV���D���7�j3���t���lo�u��ET���d�<�8�s9�?���z�e~ys�<5�kb�8��o)��bJވ9�#���2A��}Q �qE*�v���y�}�K���)N����k�N����)Ĵ����A�Dx? (�?��tE,�1�M��4�_ SN2�:	B <�M�'���Yh��2$t�|b�/i8��9w�Og�bE��� 0��;+kK1�@-���-A�f[(y����6�cD�!�M ���qkO�j��Ү�9dD�&��"	'`���C����+)�hļОC�2��9�1��􋌬�4����})��?�OM�)�J�\Z�U)˭��R��為W���\���m��zƊ����kB�\�������{�\1~'������A�X��go��>�ҳ��,Z�Y�ke�ef�݆����Z|-z}
�g�BK���@ºiG�2���4ðG#퀊�����?ބ������������;}�vG !�J��U	�R�,�l�hn�1L����":v'�N�X��E4i잮lh��4G�[��G��͓�W8�{l�e=ag�(�Ps��FOa͹�E%,��X�!��v�k}Wl�ۤ'317�Kl�3껓��S��@��*�d������SD��|���T�c̢uL�(�4��;��9� 5"��i���Fc�Ӳ��ޛ{u�wiS=.��Z�!c�}5v/����sm��a�v3�땋
�am�����<�ko��Y���M㯎��J�����x��#n�$!�2!hRVg!Skɜ����=���*�����`(t�	Cխ8$�?^�rO����rk��]�<�kR�\y�wl�E��]wa��� kK��Et��5�[ܴ��Չfz٪�b6+�ǲgۙMI���9蓼#'���s�q�SX��c+:���`q��K��^��Bdh,�D�N|�]�\RE�Q�s���e�טIC��3�=ɯ��(t�4�sH�&R���t"�3E_�	`�jk)Ô̎7"�E�N��Y�8ƒ>��L؊���IIf��-�w�zS� ��dٗZ�\�s��τ��958���P!B]}�gZVh�=�X�F�V�ygh�̽��Q���b�\�m#_Cj�}_{� ��cX༸䞭U�G��/m��#�W�m;��5��PR�zx-W�ݵvr�L�&_��O]��U^#)ٕP 	�ǩw��� �e��;�w�[���֬��,m$p�6���q���h�s�L��㕂�(��LdoCj]ğN��)�O�MtϢѓi���l�uA��?��fF��ѵ.�_ H�RraP�Q)�2cC,�kYt�M�,�( ����0��a�xş�pm>R�sZ�ɜ&}z�morNP�4��0Z�_$�ݿ�G�����d��ryj/�3�%��M���G'���.���q򭡯 E`-/1�(zC~��o�U��B*k��tY+�Y��9�k�Ψ�@���G��!���o8\�:�.���m�x��dW�{l�S�g�г����r�g2�����.kF��]i������f���#�D��o�Z�cxE��WB����~�?Wm�`Y�E�~^�4�*� �},̉�'q�Qǌ��{�K��B���#���Ҋ�h���A������x4_������=�1��0)�N���,�H~�&��,ġZ����qs?vu���Q� �����p�##0�d�
����eP�X��l�U)�9����Շ4Y��b��o��X�/�Ek8 �; �Pn`�l߶U��v0Č�ر�x2u�v����_ 9�kĎjA궣,g��u�&��e��"���O�=A�M�Z�A�U�QvHb6`��)����g�P� ���(�;f�<(./-^P��I���3AW�X���wOo���]��ڴy_�A����B�׏�\�!	���I�%;*8TZm���u��7����Q�G|�3��0"	�n�`��`���UR mI��@����P�x-�e��7m�zw����Y�]:���LM|z����{�1uY��iԤ����:�!Gj�ը��z"�)��.�t�_:uI���ԅ�0l�^��!��5Y���YH���;� U,�T�D<0�ktOȭ0 ��nʓtIC'����y	���IX�|�J)���0]�,�a�'����7@�}�e��wX���6DR_���(�z$d�o
+��Q)];JfxNn��La�F��r舁NK�1l���K^3Av��B/\��T%����c�΢1��qoФ��d ǒ���2�*�0ЕAOˮ�������|����٘�?���54�N`�U���	���X�[��N�eC6�N�����s�3��ttNja�IWW5�JO�U�pHR5d�In/�	��Y�O�H��*�w3�Æ}B���'�3ҹ���b��>L���>D�b�_?���׬��JF�T���լ���AcΩ<�ohH�a�q;��ݟŔ�4�b5��V�I��X����Gh��10��?��k�A�`�Ꮱ#�tӫ�̚�g��S�>��6E��l��DSv$Ģ�d���P�x��m�E�R |�B8k�>1��p����X���'YѨ�9&?�\U���/��G�#>'}����*���7���,����:�	>�T������J�������h��nkq�GNn���~��H�� �j%�Gn��W��Ȫ�� פ{�7F6ed4�N��Y/ɛ}*��}���K��R_Ei�ru�Z�x,�]Oy*���2�uPץt�s_¿�V���cB�����xڢ�����o�Q�._{H�j7���xE�1�K��Fj�Q�M�� ����D�ЯwhV��I�1S���i#�� �HJ�����_�����Uڑ����v7��78��3�Y(3���7�yqG�8C?�ڥs9FP��ؘM�`!]��{��b"F1ts�l��g���@usң�F��o�EO�1"�݉�	��t��� rB��5�/Pw;�����M��x-̏
� I��@��?���~|� =h�i5'�A}-I�Q[���g�*�!?�=鏁/m"�8�˹�{y�Ë��B&3��7f�&u�\ ��T�{�I�- D�ܥ��B������:w�� ���U)��sS5�],ꅃvq騄�!���ݻ�I�Ɔ��Z@@�.x�Υ����;<��)ƭsE,+�xТ�}���G*��I��׸�?�aC�Ǎ��aR���Z�]�ރ�]� g�y��X	 y�?&�D^��d?⁂�H�߃���)�K-�Wτ|p�-�#:�D�Z�����mW�"���5�|��-O6�1\-�-(q���x4��7.�
ߊ:�;�������"�ܑ\�K�S�@���W�"�ݛ�̉��ƣ)>�}dE
�G5�����}	}�+C_:��j��<S�@��N����L��.�P�)�Md/',��bÝ��>�20ՆA��٣xT�����Iﶝ,�Y����!{�/��h#M��~K�_E�nk���~�%�/�#�#�amf����y�4�\�A�,�E�W婢0��������V�*g����b3��(���=���,m�9T��j�b���]�F�j6�a��Қ`��80�6�.��zץ�!� �1yq�dM�k�����zz�	@���Zm��ZjkY�ϱ�)/ݦWcՑ��i���U��˶ŘΧ�w|2<� ��+�+��>���-�4E���}̜\�% �1��4�ω���KR�8<�')��'p�TY(*��^w�o���1W�P'4�1}O�m�H<��`��^r��Ρ�Lr����D�^<��gU�6�S�����쌱�5K���e�l����I��0M����TՆ>��G�-���_Hmw�rTV5�Z�����3�^�&�n
�=ظ�I@���J� <F��3��n�)���[mC�>��*�{�S�E��Զ~���r��R6k̖o�����o�WTJ��[_������1R\7��b-�m5�i�|����8ý$�PHjӦ ��ѓRƬ�#�w��]�<���X3��N�������皷�Y4�͢;��{�£�֝��ҟZ��q["�ug��F0�s2���H'�AԠ�9��2`#�UՇ�P^Т�G���琿`��</�=1y��pv�G��Ca�C�6Oox�I@2�C�c���Kةbp�\��Zs�^����J<+�k�7/�G��V��.2�z����]t���6y~�<}K*Lt�j�7���	a-=lKةIxM���Ǝ��fWv\����vw�1�_<;���D�Y?>���3-��2j$n)~8�nxஒ�%5��6~2�-M7�_➬"�)�� �������,B)酲5�nR~��66���/�h���y�h�e>��r�w���Z����zHAv��.�O'�2�p������v&��bJ��?Z/o��.�@���\zn���*� 
�3E�f4����9���(��pa��Z+�,�ږ@�#��	�������	e���mз"��OU8;ˌEB��z��t���QhZ�I���0�uxz<t��<l��a���Z}�dt6ì�M?��|���0�C�)(�9֘(�ˌ�!��<��#��Z��%$���N_��(��cq�L��v��=������U{��M��_��7*�\[�s���*��#x�
��gQ�L:L�l�0z�毾���=�nR�&��C� +I� IiRܐ?!�o ��9���X�K�Pkf����hз�D_+���?��7n7��Y3��Y��`��u|bF�t��FkT���Kt?q���(���8��t��Y���H ���ƀj�0}��B���I��*�t�����ߏƟ=�ȶe��������V.��N�+�I�@!?g۟n��À�_ ^�� ������KJ�p���{<{�w�2LČ)C^�O�yu����gH����aCJD���Y/²�Y�t@�쟴��ͥ]I[���^��l[8�U�X�=�'Jy�W7SB���a�V����i(�g*w�_Qy�&g�x��g7�4�����N�R��|��W�	@5W���@7�4'�L�d�$5�n�sr�+"���U����'�l�M�O��妪���o��HDO�ēdk�ϩ3�^����r �V��h�۵���2gJI�#���,�`I�(XPE�)뢘���^ � ���H�Z�0
�*E�tr *�?�P%-3+o�t�^��K�c�s%~i��Rc�9�#�=�Am���]��F'f������,U��Z����+��?�������u�I�����ʆ��Z}�멡�2��w�\���q9�d<>�]8��N����4�)�u���wf�V�e�ݵ���8H�d���t�ypd�-Hh�z#�%pi1^z�9]�_�~/T�̕͠�f��A����n�x���!����'Tu��a򕄿�=t�I�$͏ڽ7�?��{�骗i�c��%��=	�_!:cY�h־�:����|1�RaSA������\E�����q��=��!AO�!6��\!�_z���ŝ�Nj���q�%w�r6�����3N�"�R��;MK_��1�|A}KttZ�5v�
0D��s�e��*87e�����?�����`m�6�%���c�8杘�2+~+�e}�������0⸧цZ_��r��V��!=�O9机��g��/�������������طo��CV�m����+Ȅ�D'�/'�o�|VL�~,�&υswv���ǥ�X��u�}���l����̶��I����Ol�N�M�N��o���*������ �y�:�$Ǹ�>e�.K���]@��5*#��?�j4f<����o�wL>��Tq&������C+���Y��*.6E|}翕��a�yrgwu��պk	}f2�ʃt���[?�"os8p���@������K��&�o���Dmǜ� Sz��s���byjE�&*~kl�X8�3N���7䈓��@�>�q�7-�l��-E�J�R�ǎB��)��P��Gz߹s�3`�w���/�+��T��̛��G�+u���Q%����2��$ך4� o�W�ϋ�(��(EN�h&q�ۮ��z�A�!��&��8����V�D1ff���B&�9m
)sk���<�����IJ�p����e��m��3��nF�Q;���M�<%*Wbh7�t�Ѳv���#����u�K�U�Y�R�,��1+�Ę�L�4Y��P�W��H+�V5�Nt�X�x�t끧J�Y~�Srx��=�ߧ��-+����YQ&��d8�Z?�3ѥ������9�d]�N���M\;��\�`٪F0���_���fn|�K ��/�ّ�xJ"�|1aT3���(�	� ��t����}�[����<2M��^�C��6	MYD�GѢ#����Ҏ�C,��; kb�Y ���CU��˭��K.�@S�'�4|~��2,�I��d��aӿ��+f��fՓB�r�*��t��5���ƃ�������{b�� t\&��P�����uE�e�׋�$6�ǁ�qv$)�\�]��4�~�ߢ)7������j\�q�?f��Z����a��y���7K{ڐ�t� ��w:Бy��*�����՟���L��̀E����31y�A#N��H�u��GZ�*
�$ ���OT�/f�L����-;���V!hA76+�4,:|�nH~K�T��,̡�v��t;e��O�&�p ��G͡��Y�bfB-���D��#��-����;�Z���-�����ğ]s�,.6���FZ0Q��B�ۉD��m��b�l�ֲ
�b�DAS�upj5�ŨA�O:��W8�v�:�)T��=-���{`~TQu0�{�'�e1�ˊ�31�Rfy����=&�·ܵI��_:��JO�V�V���P�M�	�� �*w�(��b?d~�I�v�:L O�M�w`�OY��{�lݽ�H�^H	C;�WY�oh�#$����
�y��`��U'㙄��@>i��e���&ݯU�p.��B���s�t�@N�g�~�:�Ao �Ȓ�>�v����2�5�S5X7�ӡ$4���a̜�w�/;��Ϫir�i��D4��js;�wu`��y�D�=8��݇m[�I>������R�3a��r��n�+���B��"m�Ja�o�p�MU��a�?�g��l]9��ɋ�l���G�;Q��Ia����F#W���^�@=>��sȂ��| �~<������ӔS0j>�|=�K�m���������/w5OSHS&Q	���4C/��w���Og�ګ�G��F����Q(9C�M����� �=b��¼a�i+��k�J�<VQ���d:��|n�e0Ym�V����}�G%�����r�q��,N:%Ӕl8sH���$�3��K�+1�`����ZGk���^1�[�w~�h����t�R
C�T ���@�����7Q�0���y2~d��Qߗ�Јi�J�n��N�'A⭑W�G��潋H�(n� �ӭ��!��/'�W�X��EQS�5ꡣv�u ٘�`U�R��+,��v=ާ�7v�-��`
����p�Q��{�4���\����,��&��$%�藭Ⱅ�A3� ����;W)8���m�y�a*^[����	�������3(�R��a
��b��/Z?�[���mI?����O&�����Q�ǼN��ƙ��)b�o���8r�v�ո��D	��ma��L4x���'\���?ƒ��z�lV������OA-�n�ɃD�+er��ޘ����$��@���.�x{g<T��IU��l�D	�z �Q�*:TB�!t��13�"E��b�/�K8b�5-M}���:yBLy6�-��$V����� �f@��<V�o���������&�v�`k.Fn���śj�c�ؽUJ����q�ƩX�G�1��)]��Zt�8��3L�~qpF��$'�������(�]u��z�r������5�*ǳ�¢�'mlP� �ݦ���h*RmG��C�$�N�lO�tk��U�J�jO�lA;���B��L$�x��('<Vi�M��M��O�!ꡛV�G��`u3��0�:m,�vӻ"9�E\=T�Cڣm�F�?�r��`,X�y�r3�H�ـ�,p�-�+
�Fz�UqnY��B�����4����J~Se��Vo"E˲h�rQ�g���O��$�c���R�(n����Eh����)�V(��.���
��H����2��ѕ}�\	�EThűm��thΐ|o�c!�
��௞ �-#��r�m��%'��=L�
j*_�
���j�qy��3�0*1	�BHxa��b1�*=�\��t��ǤJfZ��x��N��l�lى�Nb�+��UN�Q6����nQ�ڭ�g��/�3��۴,B���Q�t�0wU�'Og]�	{p���}<�U��1s`U�j=�� ���<f�a���1����$�GH�M ��Oƣ#�����t�:$^��������w��n����,���8�jk2YtU;��{�3��ו�Q�d����RhʍP���ٚ"q��&�c�"*�DE�;	Sh��o��T�� ��@��?zr��C��\�8�Rha��a�8U'8q�0�z�$����b�<�(��~�`���)%���U,}�����wL#�V6gp�/3��{�p��u��6+��5��m��ى��/�s���\�ݣ��Y�+86L��K\���#�Ast��$r�u�����f�.D�+�����]R\�*��@�(�����/Ŋ8�R���QW.ci�hS�
Ԁ���q�-z�����L�'&��p�������
����`�K���ԑ�<�"�*�z%�����"��&W"Qm�h(��,g�z�_���J�����F�{6R��!_<y<�~�1u�����O,��=��E�}�5�(����x�� ��0{�9�x<�S�
|���E���M+�OA���T��y��B��mNUo���>��������UU�q�#kv��Քu&��kH��������0N�:K�Q������٘���C�)�_�w�~�`�8�cV��ߴp4]ڊ�tI��Y��A|
/k���mVĜyͬu��Z{��>��=i
B<���'�=)T^�ov�sýx9�c:gMX˜=�b�I?JI��RN8N��.�5��@���+�N67��	���6d1��(V��K�6R4�NߢqYwn�M�T�����1�gė��XGTf1�n�Jo(�+'�u�ԧO�5^��>��r�� |�j�j����}O�*Ȇ?+�t���-�>B�\;g���Y턩�6������=�eYod������ې>�
#�̘a���K/��b�<�]����{����MD�>�OP���;�����!}w�=�ʍf�������A��*�eX�2|���7P��B.����;Jt�b��'���G7/J��|K����U;���};��@][�N����$�>E�B�x0-6(Fsw��6���8��s:�n�Lph��Z?L؂���;z$�mL���w�C������>�YX�����U\��j5RQUg���$h��5u��=��͐1^��!��iU�F[�&��Oܒ���uvOzD�k>z������}�ߤ��G7а�i^򣐸���T$�&��3�<`'�:��Kf����L�g'�Y���lS�� ��JU#0
p���"ܟ�>������zB7�FĎ���u%�r��M|����h�`/�o�sp
Pp_�����D��9��~u�G���P�K�_%�����O�����v��tS��jZu�V�Z�H���2A"�~�Iy�)Q�4�[��^�j������a��a�y̗�ֳ����O��~z��h�q��pV��k�s!]z�w�
��&~�U�Q���Z~o��J��ݿ��&�s&1od�!i�'IẸ}�6k׌ҋ����V[��0��yzX����:�,'��5q����?�ܵ&����_.� ����u��n�yH�X%M{G�ղ��qn_��06��)�Z�J �~��*��I@�RH��u%<�?�Dt?WM3>傃��є�F�|h��Q����Vs{�w�[\>��{��<��^�z��ce�8R?�����ҙ�Y%�<�W��No��h�t՘�*�'�J����]���pĨ���&��g^٤ ��ۡB�v��*�L��T\�����Y��L.c�y�0��m�x{��u�*c��VD�$'b�r�p:$��=h���|!3N8��b�TSZ�vZGm�f����L�4�h�셲0Ah�õ)��khFg���B/H��)�t���>���8z|ܦ�Z�7��C���<C�$v�ߞ.���V�F����$rU�S���U5}���u|��3���,���צ�u�顦�$H�����K��5O��������I�RD�b�J�6:��C+{�j�Bd6>���4<�����c:��푝�U�=۾��r�Wg��*�@$	�>���@cR�Y��������v�EFTUǃ�rU݄���*��W["�f�W�Q�'���	�{m9m��7\*#Q69���������&ã���/�-M���� ��m*�A�ڏ��0�;|��'E����Ɯ��W^�cbm<=��u�BR5�@fo�y�[���$�� 4$ /��dT%���E�)�\&4���1�Tqf�q&�� ��^ܟC�ȸqn�\Ĵ	�کd?�c6N����K���TG��zQ��C=�s��F��wJ��m��}�{Hk�ַ8-TQ�l�kyU��O9.�Ǯ2����,��ꊍ}�+)�'��e���d�A��L+XP�F��U��\��l�=��Æ�qK(�^6U��̍r��-i�t����_s�U8}�sZ�*H�8B&��|�#�q��@�7#��GKRd4"ȋ*H-�7�$"~��g>�Zȅ	;>��x4�#��4�	��q:	��;��x�������!�]�4���N�[*C�]9��x�M��ޞ�-桱ǂ� �1�B�c��U.���h�[��-lsϺN��\���M�������
���29���6yBAaC��1�xT�,��*��ûe����������d���/�P�"JA6� �j+�Kp8TL���ۤIC���f�v�����	��_<v0w��@hx���\6��LI �i�?��4�@�nrfe��B�j�N��A������Q���H���:�$��,8WN�Qҹ�b��o�\��W�c�pm������b��C�+�K��h�l�]�F���(DH�<��O"[g�=5�G=���s&&�o|%l�����I�c�'zv́ �����92��G��R��-M;�0t�n��b�������9.v�1���O6�UP���pgV�6�L�따�|,K� Ԁ�>�\oK��	e8-7����n����2<'�) '�<9Jb5��y�pi���x��~@�77l��K|t�;���{tOЯJ�����~�p�	���/JM��Ul
x� �"�zN���a�sM-��bK��h��g�M�Vp�Uh)�8"��m�����[�/��:�U0͜���n�c�L��Ϥq�����^�����w���K Ic�����p�)2���#�Mb:fT_�!g<	$�riF����1q�&𧅾7R֜�g�<�Mf��b�i�
�����~����X2�6:Tu�=T�N�wS�-�x������2ѷ�:ܞ�}�Y�q�f!檕�����|��qmW�=7��@c�
�����ֆfWB���ԶF�����q������`�~��N�y�r*�Y�kZ��4<��T���Y�@ x��&E�lSo���;��O������okN��^��X��6����	��~h+�r�@�!8�h-�c?:�|�|e�fDxK��RC��k��WqM�ÿ���V��ʟ�T�B\G�	i�y"`4�.����.���(��/��z�Ϩ�f�]V�0:{��ו�o����L5#D"h���1�>��"�s�N��rD9}�� ��[n����7q��� ̀-��O{�����5��7� �FP@&/޳_3F@`�[	��;�)�e	�Qs�V:?�1����A-�¤�۠���z9k�
��|����VVX�m�����H��~��DZL���Fjy@1#�/(WO�iy���@��*Qtm;Uե���u�9�N���F��y�ҹ�I�q|'��B*�%�#a1c�/�o'Py�9�G ^��l�(Vf������~e�+��(Ծ!�C��{��QUb�Qs�T�o<�Q�څ.�uU�K�?L̫.���A�	L��"����Ѵ;��B���%IČ 9k������E4ѵ�k��9{�a�5�.���tS��8�[ש}���8��� ��6�9#�^ߋS��8gd�@������2uLT��R��D�S�s�˄$�4?�f���#��B�7&>�|�X�n|�iĥ�[�y~��WEɺo�Z)c��q-T�;��-7H*�@�~2449ܬ0��O�m��4@0��E.�O9���Ԗ���>���)�z�B��YUb��ڢ����&�M��$�~�	Nd=t8�vPNB�8859ˤ�6������Ȗ�Q}ƄI�\��4^}�~ʜg�Q-��Pw���=+T�D�e��	մt��d�YG�;��N
�=v+]���@t�t����G	�K����I��4\����d-pH9��`�ϔA��j��E���Q�EtDtW9f=����w�P��8]U޹���ˇ�q�+���zb�_!b�~������{��ԧ��<�
y�����?r��ɚ�/5'��d7��'�V'�����RZgp��y}^��T�A�o�	>`wqG�\�S�B��=M�
���dG�.��o���9��A�y�!�"�Ni�h��
��v���oz��?�%x�?��;��3i$�0Q�É�����P���^ܰy�i�*E�Y��w_Zd��a�n漀�J���s�l�S�nZ܅�O:u������3�����Lx
��G|Q���p܏�"�nm �^��|�=+�o�����w,�c���1�g���kR�ʅ|��&�V����cp��e�E����<f��k��[%@C����`�8>���a��g2<��QZ�
��j�m�������*h΢�.������':&
��i�<�h�1	9lXQ�q=<-�y=��p����/[.�8�%"J�+7�Z+�9ٰn߹K�J��-��ZIk���G��)`ͩ�m-)�7��#�h{ļ����a'��r�I��>�ʜ:��M����K+�J�avSW�F�y�
�����&�FI����9�,_�dR/�a,�ٜǯ�	�j������H� ���s� N�ű5")���������	7���v*\(�
�g=Ws�x1�P��8�7���C0\va]���l��w�4&df��C���@i�}�a�lYS?G�,Q)������v���e^C,#>7Ru��ZW�vWa�iRʤRubxgy��j�A6��G���&�P<I�"Xfh_�#�����<$*$�6I�}��y��U(��܉���˖'��d�X��=RPw����%�?�ʞJA�^��9wx�aIY�x�j�e��W���3����MA���J�)����5�h꣒f����1$��:!I4���6C֢�[����UҀ t@Zp�R]K�D���)����VEa�:]�/``����0m]��$o�
p9Ǉ�!"	:].�KB~~O>䌮W"�fZ��B�	/�5��<d
���h8�6��@"S���<�.�&p��>����=�um��%n�kJ�����:e"/��Y��04���g��N����3Rͤ��UQ��V#e�Z�W7��Ӂ09�RĹ�"�;�t��vkd=��=�[�H�	�CNOi/]��"����$�ޥ��Z_Z�flq��no��N<��<�X���y{(>�1Ìy�ഹ�4v@��d̪�.aG�ql�iM�ޒ��놰��^�/�����\Z�������x�������%}�h�d���90��	;�paZ�K���MA)Ã���1\li}��+O4����PV��(6����Ix��ٶ1��,L�E4�a���$��}�۠��H����5�R�Oz�/a�X���y)����w͉a� �$h�$7Y����6�6?��W���I�����bQR����QEݕ J���Kp%�ey�+_�{\�{�9��4���XO3e9�K-e�m��2��v���	B+�%���.L���,9��JQւ���-&ό۽�Y>���6�Г���kWȴ:�������IV���ᵴT��K��ِ��_0%?��]�{�4j�p���_����R]��j�yE��t�R�yb��e����ڤԱ`N�1B�bu�5�>����ȿ;��W�QY����Wf��x�0z��s��D�{N՘d�E��U{� Yhu��΅<�u��v�R�(G��N�$j��5���Bِ�CKh�>L}��]��biDuR���>�]�G(32�����F)�>��kE���q+��.���X�1,"}�&���A3ԫ��W���ύ��=[��ݚ���Ur�#�F~������1�H%n�EÛ㿱D�su��ɢ����!��J�]Ge�.F{"i�W�m��|[�<<ʬ�vID=A�>�%u(Jl��o�X� 9:D�An��hjҽV�\�˿�8�VuLs�w�dz�DP�%(��y����,v�'���c���wS��y^�+F�Ğ��ؐ�N���,�.�CI0a�4�"ʼ=���q6�K�"�P�1]�7`�z D��>v"aC���`ӧ���m/PM3��>�MQ(ňe��Z��5`�@��fw�\����h{;�D�v��6� �x���"x�	?�HO ��<1��y�`@s�,���5�s�]�v����CB�-��?�^_�A�t���J&2l8س�wf}U�(hNQ�ED ���t��f�[�<�Yb��OoֵV
�k���0I�4�s��vձ��Vȹa��-�j���M��!]#��D��+v�~��v�v��Nicf��#R���HyTr�B� &���6�}�-�ٴ>��Dڳ�~�2�0M� ��s����Ti�K�H)k-E"��i�7��,�,�X� /��4�R�Y����h%��v}����Y3U(�3�����q'��f�]h_�1,�� ��}a�(�@	�*�!9�嶻I!���f��U�>M�F% $w�6�}�n�IݝFW��P��1�۫� ?:��q�d%�����O�!�p�G��%@0�̓�W������22ݭ�ɠ?�S|�Q���Kt� *�JZ`)�XM�:$�5��!�z�7'~�LX7,8L������몵9�@4�n~J^�Qx������G������ͩS�d��JG��#$�����2M��#(��8*`,�]v���gs�GB����Эm�p�J>���v�R��T3͋��U q�+��&�25g�J����O+�����[�{�����ͭ��b���F�״⊤5&���:G��X��R�I�;�yq���W���!�C��4�i	3P�9��6�|�2���J!�������'�Hn��a
S���PWP����SDv|�~ӊ���J#\N6'�a��)�S/m+gB�c���R��&R�/k��ױ���΍M�i�x��
ϋ������F��7�s"�C/x�ݦq�!��\=��On""��t��Y//��~ᆗ��/NT.;ER!�c�L�u7�YR��歩�w�`��a�U�~q�y~c�+����c�k���]%2�������5�<�y�-�{X��	����ˇ�ߦ9g�|)Rt����d.�	�-q�g>����`��tJ|��4���e�:����1�s�WН�b�U��&�
{�3ٰ��`k�%3����u�ͪ��r� =��q�v�).E*`(�k�K}�qB����\>e-���x��1"<Yg�����L�f���oO$�V=f�T���>Y�Ǣش$ �Z���,�p�|Y|Kj�_��n�@C���7��	��w~���c��ڠ�����cO�*�#d�8��X���4��nso.!z����Ј3����!>�P�zu���a�,U��1�a�P�b*9����8����g��n�)���;"��H[�Z�����i>tߜ��?n�+��֙�	�h�u��^��n ��v�`VS����^4���W��� �;h����<H�ߣ���<�s/[������z���vh�	�g9<���H�+r�Z��%/g,9.������8�1;cl|��[�y�H)x�Sl�񒵳�`���V�׋7~���{�\��Dn��}6ā�2N�%Bðd>�\�.٤X��hձ�t0	���+7a����.��P��M�,�]º�1��भ�f�(������N���c��/U
��!���).5@���m�(HE}��Y<K�Ú ؊�9���Z�l�>�K i�z��v8�ewl�盉��c��|N�D���u/���1�W����
�+^/���F[��4R��%	6:+���_��F�5f%� 6j`����;N�ҧ��F�IO�"��j��	�{O�U�~~Z<��$-�!^X��:��|��E�Z�ɿ��ZKUkI�;��b�p8�,U>�պ���/��**T.xe�r�JJUm���E��C�~�&�:L}#���t^V�Ӭv�덙��qz*��I
4�b(�.���v��]���4'0�ҧ�Q�#6��"��2�R�	xf�����*�6�Wt:��wm�XPGQ�ﴕ#&U�ڤ-�;ە�x�G�@�+E����p��\J!��#�o���6
�X�	Ϩ�*������H�d}�$���[-)J��˪K�7�uGؚ��^K+*�9�j%{k����9.��?��ꅅ:t��[I��9a�G]ĉc�^��H�����8`�D�����<���"N16)�꾿!a�,L��5Af�<�z�.ucAs�q8�I�N�l=Ց�~蝌���GX~�L�Ê#C5)U-�F�;�>�ƖT�vj�꓅^���E�C�������c����>������|�e��3��ieǁ{�(|��kjǯp�j�m2)G���>Z��`�w�]X�$���/ku|Nb�G�y@&kO��h�g�{�>� ��}�h��|_�#^�h���~���e��2�}��d��먨^��E���:�7
��}Z �3�)�Y���w2R E0�ֶb�bB�3���?�2�U?�H�9]�b��;�-��Fqt�t0�ج𿊇�CZ���}��L/�kM�?����~�:�R1�=��>g&RG@r�o�#��>��=^N��q-(ᒅ��tB����%�����3�L��r����T�W��#�L�M��y=�
�0X��K�h�c/���Q�>?�P��c"���&3Y��x"�=��%�m���	�I���U,���Zk4ET��?�rd��P^Ȏ���fB#�&���2腲���<���4��-�J�)ē�b�'�g����<��:-c�L��ꈃ9M-��u�H����e���͂uGР����{c()Qܠ����������<��o@옊���#�{�H�a�zu%����E��T��K苒?�QHW
>���t;q����R~��j#J�י�å���=� A{�`�J���JR�����2<���<�5,�b��a�B�b�IH����O�N�/TՀ��j\����9�fѝ�؏u�Y4M;U�e���y��V�5�&+�A�rm�"�o�tR�e�/�ϒ���*qˡ��N��߬$�����6�(�m�VJ���~>ie"�t�6j06|�ߜ�z]�l��Y<̃3��R
rh�ტ,��
S���T�^ZaU�y��kp�T�}� {E�8��37��P��wg6�]�qG����'�����N�hn��Z���2��W[`!�lzQ����A�i=�3�=>��$R�nt�t(��"� �I��Mn�V#op�/�\r"����.������"o���=-2�*jw[����d*zh�����ն�:(��*J��1����?��S$��iB��*��B�Y&�����g�>X�GH��,*�AL��Ty�7�7��$`Va��Pî���쥉Ő>Ζ�o-��6p�Ƴ��mE��m�JmY�n	,�kd�5ՃL�Se�|��JQߴ��d�l�Sl�fS���l����`{� �M�c-q�˦�[�q����"�1�T�ۥB���3�*��2Pls�O��,嵞j�d�zvG�#巚������"j4���wn�B
��\�K�!x'd�&�Drx�����bq-s����ϊv���]���&V��g�����?��x_��{*<��'�a�2P��
$�Ǹj���%��Y9�"W�eɫ�o�r��i��YuI!�Lǅsf������7�t2��r��$<ob,i�(2\$���$Rk�)��F����XR��<���m,�a��l�"��#�ޕ:/����©�nG��71RbW��pJs��qS{�# 7���:�0�U����T���s��Ղ�e�ќ�.����8oF��!�1��<Bj,�4�Y���5vҙ�!����dd����k�fE֬����zc���@V�;�Ba]�����mՑ�w79惎�U�B�/�{p�ԭ^|>��kg7�t	9�(��"����ӕ4a|��zp�:�-�rl�	�w��6S�K]��!>��',��7���ݳ.}�l.�Y/K��|�ߕ���m��1����0$iH;���*Y��0�؋Z��@���I�V6�!q_f����*�g���1{23��y���F�.�XT�j(�o�R�T
9h}a��wQJpO����Z"%�S���w���vwz�=[�(!�U�m{1!}��p&黗(@�}w�uM����A��!��/$�m_�����7�զ�h�F����P����y�S}jAo(':v,�ĩ/_B:�޸��~��͆d�����-�qR���G�5�V� ��'|1ON������y�������0@�B�|�*��M.n\��aJӏ�j{���e�(q ���'K[1FV��_Eu4��n���hW��6�G���d���6d�c��"��m}��%\"H�/�xp�#?��y��\K`��Q��|�	� I� H�׮�nu��Rq+s��Z��[��#��� <'q��n���lEQw�X��ŉ;�(T�díB�0�m���s�z���/+M�20��+��Eq�����?S�+zm�d(2Hڹ�,�c� )�]e7_�ok�
L[b��R>��{�Q���"jT{�8��s�Se���$6X}����Q J��Z3߲�T�c��);tfΩh�*���x�#K^w���م'.�S�K�˥C�Z�� A�N_-����w�OG*�dl���rˌ8�S�ʒ�⽨��Ϫ�W��d�"�ؓ��-&��L�V�Fw�턇V��X�ȱ�q�r������q����#�>0�8Sw��gs%q�@�\{��'w��J:K�`��w���G���C������$�2�k���`=rć�WF����S7�����m�`�K~'ԕ�`�=M}2=l���1�Qt��u,$��z��y��k%�ӎ�bE�b�/Q6���C���[+p�Y��ƏxB��K̒�z̪��<"����6�$2��0�D�Ah��a!ӱ9�|��;"��V.�>jvm�s	�Q �XnU���	�<[��+,>�D�u��m����0��YB�����6����B��9L��C�4�Y����[��kf��d�*_�����ύ�=�?sЏsÛ��K�\F�g��Q�@I�t&@yGHm�MGkbH��H�H4"$J~o�d�T��(�,`rb
�B���{��0��|���������đED��v�'I�h��JI\0�d�.ե@�QR���N��V���g�����]'I>ȭey�����D�E�$��m,��19�jnO�o�/�������jT��۴������X�Ġ�R
�I���$s��I�Rb��e�h��V�����Kƿn�]w����Ey	3g~xZ��ݖ�j�K̓��͠�����"�`J��k���p�������+�s��DleY،Rpv��y^�������kH�p��������M��>̊�T�0��EF��YV狪i�>b�Wq����jCꡓ@��D�x�.L��./vw�Q�b8Xs_4�[�p5L�fT��D>�$�{����D������J�QO� ���idsJ�?Em��a���=�|��\��>��9
�yP�s�[��܋O��ǩB��/0���7�/C�Q�c��)Kc3:���@� O��H���(e.�R���q]�n	�*!0S��?x�A?[��VyC���MwE�oa���Nr��ԥ��OD2�I�z��&U��T3e%k����Ia��v����R3�(��6�,�p3{�.!�uui61Wx����6��bh"�_԰�|�*���TfW�ڳ3�rA�h5Y]y�+U@d���)�i��8�3b�/�8�{^v��P�)E��"�~�{ΛI:�,#��� -ԦҠ41S�������8p5���N��p� u��>T��;�@��<^��HK���C���	]��]#�FC����F��b��]��N=VrZYˎw�>������ C(�.·>w�OzpK�1kC�U�pd~ick�����H�e� ����p��<5�x�v�=��y����&A�%�]�׼a\��C�a���2�H�-�D�M��MIXt��I�UcM
XbPK��8G-Ccwep+q?z��H���ͫ[b˝<�Hp��U�@Xw��P����1 0��5we���9Y</h;���Sha���7�n�oJ���J�O%�>��BD��.0���A)�H��str������Ĳ�v���$ݕ��;<:� t-8ßN�Y!�"N1E�CB߹���ѱ� P�E�3̣�W�@�T}�By�?�� �4W�[|BgLܠ�D�ִyaq�k��i��.Y��:���q���ĵ��7�T�N=��,����d���;~k�^e�
�;�o�m!�N�VGO�3ߏ��D�{�>��J�� !5�!�K&����(�ɝޝ�ճe�7ʅ�l�c�VlRiW�\�j��}[���@�6��������Ð� 7l�XC}���Ƨ�/G@`�>��=b�3�BM��,}Ä��S'&Q� ��+a�f���M�
�S]G*4���t��^K��)U{��~��t���T��EX��D�/�2¸޹O������,6Y]ݰF2�}O���MA;eٰL+@a�~�����UG��R�<N�����_%�u2��Ey���\�PY�b�ŀ_(�z�Z��P�ۨ)�z4#D�jഡ��L�����|xp'����O��%"P�lE�'o��ї������cc�!�:��V"�j��L�͠M���oi��l���� �w"b���~�]�HI��Za������d�`�p*@~7WgSbu��i���'5�JVT�@�&���6D4�:�Va��v���q��0f�� X�Z#I�P"�.��K�ȧ�1x]�% >+��⚸�\�$��uo���L:C:�����{~����~i4<��P�x��%�
���9nR��Al���ʯ�C��h�'MO~�tPѺ�����^ ^����j��+��sb��W4/�볤�wX�X���B� ��t�C����Ǘ�s���H��䉏y#Ni���������Y�	�.���u�k1���J�2o���7d_��sC-ƅ
ׂ�:ȷ�-u���V���<�.fu�#pZ1�d �L)o�p�[��
�F�{:�ɸ���J� ҘJ��`G���c��Ew�sm�Ѹ�ӽ����N�m�r�i8��d4.��~�G�P�1��	2-?���TTP=b�;>Z��"�r���e]��[��{�b1�'����;|������RG��� ��L �~���g�����5�um]���!����0|J����751E���&WA��/�I��7��Q<�f^��B&�ǀ��XH�5����f�zm�8O�)D��S���u��sd#�5�o��4��R��JZ�}�W`=����9�3
�ac׾��ٶ?*Ygid9��iH�m���x��jC �s1܁T���.�(=�@r�u�L
H�C�<N#7	����$����";l~��"��X&*�,��].ؿ��'�u.���c�`���rX;��4a�1ĩF���_1˕ow@��?���Z�����Nö4� L �Ã�rxI+2,���]f���۵[A@|�����|�qp��2.��Y��>&��L΍��	�E<#J�����.��0H>Bf'2o��W�����u?�,���tR�����x�}/\���b=�*`�_U�^ɵjIsY����Ȏ�!�rG�����{	3����$�b6Msl?7�o���	�HN�9���}@�Ĕ�'%*^3�`OU������? �w�+F��֤'��!�\Ů�IU�a�$��|�@yީ9ޖW��?>�8�'�4%Bg5��8�� ���Ն��� +[�ĝ�+�>�s���!l�^s���fRo%� 9��^y��_a����\K��Õ�KI>��#E.,v��2�:.���f*79�.ߝ ���O����K��.ɂ�����ͽ�ц%p�:�W�Z��^����ç]]��r��v��|�x(���}��8��։6W?��fK�mZ,�Q�5+g<?Y�"��r+�N� }���w^�',Fy1=�QdI�$�E���ɉӒ����������/�5�ݡɜ6`1��T�ƑuP������b)����k9���iJ�>�"�Ȁ�Ҷ��|t�`�tl�.^�d��KL|"���j8��\"Э+-����1�2)1Yq*�~�jh���~���L���;��+�v�	��	 ��λI?�v��7"�O<���:�{Z�-|S�fO_����].5?�˓�fF�@�bKe]t
 Zu�v��%2�I-�-r��'��2�Lj�XE5���V"/�V�ׁta���P ?g'[��Wo;�	E����=�e	�ˊdT�x�-�� �RL"�h�e��hg�"M������,���㸭q�F�\�B;���_tK�w�����F���B�S�� ��ȘPAYJ��������P͟6��k�.�~�`��uF3��e���Q׼��S�����R�����J=.L�����di,�T;�a�3���P|+xe�y��9�p�9 ��,�Tx����̊�� %�,&hA�~�̈s'Q��"ɾgl;\/A&I����/�h�~uܺ����"\݋��kD��O��)���'��+�c��� M?vV' e�;�*�Dx3�%[c]ڤ���>�cՐ�ī�<�{�H�Za	2����[D����ü��k�ф���D�x���S��X�y�}=����n	K?&����g���L\n�pH ��S�Ч��G�c�����N3�3�q!����#rZ�[��Z�5��U���H�E�O�a�Smr����Nw�$�9���r'�� 5��N�d��H(֍΅�SPZg�9�M.I�|'�Sm1��ȗ(���y�&��4H��@�{?�ra,�#�U֩3,-R��6�?K)��FG�>g�0"��I�,/�or�t��1�q������z�����r�ґ�9�>�k`i#-#��Ɛ��p���Z?�u'+L���c5��BB�u�5l�t�%l��u>��E���<��zH�T]u$Z����a����e��?��Kz����]a���{�L���ߧ�(���Ӵ�������	���~����meSFm6�p��Z堛n� B@!E���p��^.I_��\�<ι�a��k����J�Ւ��'�Lcp�۬jz<nJ9�����תSa������5��=���؇����m���7��D�vS�PĖfu5=N�~e�5H-�ۯ�=yh�cT2�h�����o��L�{�Y��K�YO�m�������n���?x��B�x�V��λ�@�er&�&��;.I�����X+v�6S��K���6���c� �5���c!2��$L����mYӂ#J_�������x��mf3-��-��G�M��8v��>��!�h�11 7���V��A���2���;e�� ^{kO�D�/�/��׈��� ��7|�V@*�8�^*{3YO:TCiv���G��. ��&�Q���4�qSpV}}��8�B����bv�{	�3}��𠇡�&���4��z��1@+K�(��0�t��i��X����j/�<q�ǔ�g��r��q�W6��{�(�_1� �)�ɲT���s�5�_LG��<� B�P��E��P�0�y�zQ�Wd�~ڄu�dS�`�ܱ:��p3���m:V��l�Z�Ɗ�i��i�6�����׹��l6f�<&ʸ`]�P���>��)`Xwc��vǶ�(�xͶ���>T:�gJ�L�%�Xm>l�y^�}\�1����y�W��{Gē���� /(4�U�F��Y���5i`��v�.�OpWg�>.S��.5���$�5�ӊ�4xF�Rs�-���\�����t�c����9M�ԨT����Jm�\����t����ddE�Ӹ�([��.��3�'ӳӱ��&;���z<AiZ}Y�yF�b���Y�2=B�t�FTk��|PT�W��I;���J⁏���kW�l�lb�ސ����y�g,�X�hy��5IX�K��1 =GLd���|a���o�'T��Û/�ˀ��	p�[�&S:.l���R9J��ie�hA�-�>ª�-�캋v��m7U3|̯�}�
P[9�p�?_:�g�B��,m�X�ԡ�&���MA�;��Z��3�7��r�4�݁@����s�7����+@K���Y>�[B��ߣ˹�͖�X4統e��_[����^s^>�fGs�9�)w_�s��ĆOt��rA^zR��t&
��치�3��i���9
�� ���A�/Q�p-#G3� �#Cq�����PJ�R����J���1�ՑԖ�9���b��R�i^U����m�[Ͳ>=���2�u,�e�����doH�_84J�/��@��[2�$�D��>e�BuRMW{��GՏʐ(4�� yv�m�Z!;���5�cK���O��.0�j�بۙ/NBEk3d��WQw���0v;��2y7�}�?I��5���l�c�0.�g��<�c5V��w���0���k��ޡ1�Yz���<]���5ca�l3�����3j��˺%�,EAR��d�/C�����}m���/?�����6`�7���t��)�:)e/a
��1���ؤ��KC:�nWX'p�u4��8&�	��(@��-%����v��R_������/��J<T�G��~4g�A���%�hTl�Cy��	&hG���ܖ���h`�w��YEC�FC��U��u�"y!#j��g��W�Z��4���'��V��|I�-I�%a؞�G��#�|$C�e̒Q����V3����I%LD��` 3]�o?#d�?f�$�̭�}�g��<���|�1Ҷ�U�~�vK����`x2�f�;F��Ѩj���Г���6�x7
&�FS<s�7���������*c	�D`v}IR������-�Í��n9�XBe���(O��` v����Q���y��K����w�@��B=����s�3"l��j��{�թwL1f��|#U�?��z��u��A����� �w�ij�� ��pW�"M�"#����*t�6�la�)�լ�U���� �G� 3r�������c|�*a�Fd�rA�%�����9e�I�U·���#���޵u6�g��CB5�X,�
��f�LUv(I�.97�'��xߛR~� �(�p7�4A;,��+
�|=X�dZBHI坳�3��Zj�z���⋕,�l��\��i�u���d��v��J��l>�1k���d�{
�`��=I���\�>��Y��z�����#
��Z�Pࣴ�|o�)�{���)�oV ���d�6boθJE&ࠢ0E^cd�C���1�4Z|��x�}�ء�?@e�h�������f�K^#2	D�I��.M� ��^=�'�R��M��+S6�,�N��%1C� onF/��׮w�����l��֝]k��L��X~����wC��2� .s�1����Z�F#|I�y���o֟r��/f>�'G.r�;�9S�>����3<~@�������%��6����B+#��K�E���<] K�2�Ǡ���0g�i�#a����E��Q��U%�R��Av��!��h[:$���%�&w�c$Ò���A܌�sC���^��X�4�{5}�??�Eb���Cg !��Ǟi  6�ܼ����;iݖ��P~|�GhP�l���']Q�8�~~�7��B}>ܣ�UE)x9�ǵ��j�b۞�^��_W9�fݾ��cԁ�oR�QȪ�
�u�����p����!L���-J3��A9N�z�2���.�H���7�(�b�n���o�#�%�ՠ#s�����,�+�Q�.W���l�4�E���ྖ��"��B��h*����B�ਵ���잠���䠤������]�s���o'�'��om��Η��~����M�����@��nט��W���jd�M~m���?P�q��0v�[���|����,F{���ۇ�Vm(�R���Ed�]�3�'z��
+{���{{�}n�1��l�4O ����"�z�C����׮��@�Ԕ֩�;j��U�7��j�el��"�BwY�Ah��.m�.��[��:e���)+�@��!��޴I��z&��=��r��������}.�C�MϹ��+8q�����H���TNj��E90E
��|��.��+�$Yc�z���4l1s��p����۬�4{��E��3��k(��\3�A�ad=YM��b�g��
�&���ݻ{�N*�
�tT�{J�@HO��u�v%��3���~[v����LG��zpRt41�o�� �=A�U�S�P�ŧ�$*��m��&^^tnN9�inP��ԃ�����y��7�^e�F��'FAl^��T���ؼ;r�R�A��>��|!(��:�$ogq[a_r�i�&�gj���^H����3k$�$�jT>6ɿo�GK>0a:�f��^JNN��f�
�mÈ���\ϼ_�3��W?$OX�F�`���F`���tb���/�o��6Xc����F,��T��T��!�W��,꿀I7��k!:�,�����,�6�s�` S�;ָ�̖|6�]qI�_m�Nx[�ΉV�~��E��-��{H�]���<��f�5�tP�� ]t�Ͷ���uUHX�o'�<��g�9ڣJ����"٠!�5
�U\��s���$[WA�=�:��TH��������&��-���c��J]5��>�0���C�z�HLu�Ee�8��IKv�`��T��✌	��tZ bF�	��ަ��$P-8uLO��������7J�K��w1���,�ᓅ�}ßG�s*���{��F�+�>���/��I"��F5vE�g��	������Q��q�(�{S�����-��7��ӢӅ���O=�х�E������������e��س�=v�`��.*��RR9�~΋�u��9J"�<���Du�D��oqk\K�Y�pd��<qS�k`�S�Ơa�0`�h��Ʌ+���?���Ѵ=]zcj�:&|�(�Z;����M�>C<C�!�����Ox��,�7O�RV�c��j03����O4,��V� $@�B�tG�� ���R��Оa�+�a�9Z�Ǹh�Ue�Y��m'8.���
�st2)�6;�t��#�IAI�i��ox	��zÍ"�nz�o4(�Iw@��We�LA/щ��&%�h�Cn��������������?�[y��Z!4+��ޟ�tz�e� {�FB��el¥�	��0�����:�s���:+�w������|��VV�&e��� ��&��%?��k=aD=*��o�.���mΦe��u)7 �@��s[�]6��G��V�*�/<Ȗ� rf4�� �G���+.C�ƫ}�}��7'U剩g�ַK>B�mπ�:��`6CYe��8I�;���P����sq�`�˭�ǘ����G�������lB{|�3Q*�>�#d!��Ҹ��q�Z���P�O�.�����ɴ�3�6(��&љ�G�"�a��7�Ő�kƷL׮|���\����=�جR��T�󽖊��	x�.p���+7j�^@���Gq�T�=&ik7y�;�G>@���,/�0�� �	Zǯ�ǭ>�˫5$ǿҔd~���9){�Ig�Y���NT�S
z�Ϭ@r����v�TJȝ������I�O����%�:��#_o���D�n�ch����*�e,dd�!�uO%$Tʚ{~��X����x[�"�V�4�#i�vc	��ƀ�:E9�B�n���-���/!���8Z��E4y�$��rZ�ɏ��c�57�YhS/a���9��9\o���aC�UC@��>H��,��ש�"f�P�gYS��<�����D^�Ks̊Rj�q�g����	�6(�]�!�]-�_{6�W5���bC]l�G�P�����s΅2�'yr��6�� !�=>��<���4VB��
1?����X(�Uʄ޹��%Ab9T�Z�.��ww�K����Hp��S٦�u=�]�� �ubV���&�л�މ�È�R�h�� �Z��i����-�����F>���a�+�i�K�p�����V���TW������?W���k��hl�ꔻ����D�D�,ްr��뷐ii���p>I�J���/2�|��A2w�V�F��'���]4��nwp�iT�+��צ�(��:�����2d���,&�UO8�����)�8zT�
�KC��Rz�z\�D���NZ�?�,�h��V�^Vs ]��v��k6�ef�V��CH�	��͏����������(|�� fR�{�Az���EvAp��k�?!:�kn��5(*h��[!'
����M|��%���*&z#�C�զiS�^� ��o�X��ZH���б�R����Tα�G�6����~ޕ;�&�t���)
��B��|�z4��+Y�쳅6�*�����Rş�)k��Zv��X)"�l#�Sn+�_j��7�E�l���m�Ｙ��!�.w�!� ��TN���&�z�x�-�_�D0�My?kP�x��������5��h�K4�m�x'��ֻ��F2�`�c��6!���o�$:�ms��e�1�o$rm@��q\��2�vY�� ��G�.��Ч�h@��r�>-(2���� 1�7�A_�T���A1�P�@���:
��~��xn=��阈|R������<J�S<��}����#����dh���0q��o\撈�)�­�^�AĴ!�il����0D��uY���.LX *W�o۲%i %�M`��?^���}���C��@�BɤPB����b�Q�x*a3��jp�S��c�c6����2��<~���Q|�A�ӜAO�۞Ʃ��ߴ�P{��iǗθ�p3��}��ƕG;!���a��k�o�:�O��`G���b]}�S�,�:tO�wrFSn�N��*�Z5 �c�3f����%@A���w3��h!o�
��?'m�	9���ד�+���rM�?�k%p\sz�x� p��,jGu��V(�e�]���6�"���Qj����?6��UN��#�T���Y�X���?x�������;�����2?�����)#����0����\���==�ĉ��"�%���w�w��ܖU��,����=�oz�Q��5V�2,��W�K�tP���w�A��a���w��P�S9̻�ձJ�	}��q!rD�Ĵ�~x+����ƺ蝩i;H��CImyr���/H��ʹ���G8�J�$��Z��0�:4��m'��|�ǟm��;��:$���t�y�q �ـ���Qn�����˾���n�#�]�%4�r�9���4�Εs�MnX�2����D���~��������y�_x�G��\�:b��5.�Z�@~&˟ ���Z��k�a��F�w��@Hf��A�3�X����8�63��yzT<</�^'۪�ю�X`��%8�Den�Y�n�}�����Ӷ��(?� ǳЛT���l�+��G����� 4�������u
s[� ��>3 �В�"�<��~/�9��)�
�tt�3���R����_���׋ۼ�H�c���N���+�l�P�6�m	6�l�2������3o�i�+�z�<�x���C�:��VLס�`�ز���^�#��/��VF�~�F��*q>$d���_}A�I��$�Ω;�V{,y>-ҕ^B�0�N�k�7�����",am��!�����sZ��L���{X���s�����@C�#!S��/���V����N�v��$�N� d�Q˿慝cT� :.}�f�;v�iI�����˾����fPM7�Q*I?�
:�dy�qw���;�V₴䴛z���٣�/���z]W?uRX_ �r�6m(JG;^��1��[��O~0ҖB�����.q"��a�\P�4|���6@km��v��<�lb?H�s1`�*c)�cu�՛"��n&�o�1N,�)��d�SPI�8���u�OkǶz�������V"�\N�'+.�q}\���Y�ii��a�M���1r�\�d8Q��.;
%l��-D��ȉ^�Z;9�����s���Õ��/·�>o�%�%��:�mk��_߮���
LE�;��Ź0�W\�=W��2+bB	FgW�|�	dQ_�6<�Fî��!g�o��8�Q6�V�Ϡ>�ʁ�O���z:<34*��3-���B>X���0���A'����]��/�T��/9���0�V�\��\8�2������r>���ޭ�QND}0�{6 ��>�#�e���B��N~7C$Fܚ|���\�6���@̧Ԙ:w�����)��Ed�V�f�hY�j��z��n�-��� 1賞S@�)6�`P2���T���S:�,�/'y��>�'_=+"v��G�1�L�h���)!��令�3�(FB�.������B�A)C�bX����K��]�JL�o'�����I8g��С��K�2(�|�q��$���n�f�N8s�O�)F�QX,���Q�ԚAB���$ǌ?w݆�(8W��1C��5w���Q����s���=��Ɣ�I�I�!YLǩ�Y"ݵį ��W#ĸ�2���<t��ry;�T�Nۗ9�|o��T���B}�ߓ7[��V��dw1e	M��lk���0��uO�T^�� ڼg66 ��]2)e�΢���Olh	�����Xl�Q�f��iJHN�j�o�� >�B'zBۣhr/�d*�w\���qz���7�$�>m��?�T!������T�p�r�����[��q-��H$��4� �ۘ
͵�����?�%/�&��b�u�B~�t����Y�+&�1y�n):�.v��)S�4K��Ɣ�����@�����\��	����z���z�t�m�����Lc��}���k�~��VDA��e�t3+�#A�t:�xx��]N��[48�XQ#�D|dGa\\� Nˠ��Q�.���j�A����7�>P��dJ%�������Z���"��7�������b��r��ΑT�kZ<M��z(eN��M��Sl�U熁�Q�OѰ�H�9%�(r`,|4���>���"�4�Y��|�~��Ȭ0�މ�r��7�rϋ��-2y�26�5��b��k�cw%Q�� e���S���k�7(q}��͎�m�:�i�J4�|�n�LIE�4,h��W2И񛈣�1�qؙ�q��Q�����*2�sH��f������!^���7�ץK�����@շ�|�/aK�rڠ�B/��B��>��.�E�Z�ߗ��!n���I,����Z��t]����s��~A�,q�M ��2����.R��ϼ�:��Q�S�e�/TJ�Ǜo�o�d���L��f��_��m�J8����Ϧ8P"�z.�]RP"^��k�c�3Q��&�QD�g��o�]�o���i(�
t�������ö�u�)�E$���Z��AĹ�4!����&9���V�%���g�8�h�]��3F�5� ������ޔu:�%��%�>�cSf�0y��u(��dT�x�M�q%�ѫ�|��(����A�A?�֎I$�<>���M�
N�i�(/�wJc��s�*�9��uD^���2>��+_��k����0�� ���u��u��ӳ;��4Z��}�*��"�����m��{�e�u�Y��!ɑ��ʿ+X���#�lV���F�`��3��p�ܔ���l�&�Y��6� w}�K�%��/���+?E&��d�LV�
M�I-z�;A��$]��w�G�����6D�_�!�����g��W@������I����ȭ�N�GP!q���|p�7I���>�DrX�����R/�K\ҏ>`M :�� ����B����Q[؍��y�����e�5d) ,�L��� �N���m��Mj)�_E�o^J��&i�p��"����q��+��,o�g�ˆ�L�ٻ|pJפ˯d�x*���T�0Z���z���SܿKI��_nV�L��R��x�}L�D��2��T�%�I����P����j���L~ 0�)Wܬ��t��	�������1[z/��`,{���f��7B��m���!��I��5/'^��E��BRZ�n���єdkӇ=�<���}xiC7�3@L��k#�3�4�ƨS.ͻ}p%��8�ߘ��P�j�^�ܾ�ǯi�7H7�s���A�r�.!����7�/ݏ��^e�˻��1�5h~��+ �^���z�!
ܾKob"�OT2���8���U�+x�:�d����R}�����-3���޼阍�#�/��YN}���X�e�"�C�e�|F)�r�u��;>FY))aZ�
΍�0U?���=r�5���`I��pC�A�o�'s(G��+!�SM���}k~j�!c�!��].T�_0��P���8��~^FG'i&g��@HKX��*�֡�n����[�,6�v/7�����)"��������,f=���7ƂI�%I�q�(o�<��T�H�)ߞ���%�t��uXg�m7X�d�~�P�_�*�Y�>��l��	5ޜt\;aS��c�Ref�tf��4���{ ��;T\�^5�R���9�z�}ex�k71��\�7^P.)�u�r��[NXN�0�*��B���A�]�P�6���c��w>=ٔ��h���rP4�Ve�� NWz�B�q�K ������ř���z���k� 8^x��P*N��97���?��c(�Q���_�Z: �=Z]��es;��B������ k�P&P��|��R�'���s����F$�V���1sL�V��5�0CiZwّ6��*�È�z���>�|G-�#����0�s������QGy!��P�F�fmR,U��E�n ��Hr1��U0z�9ɡ-ث֘��q� c�m����?i ������L(:�������f53�P��9m�zp9�������� ��������:;PW�ϝ/���,d�,�Щ���LkjQ;�W���2�Ǫq6�z8㠒��+&H�������[}ߍ��gխ/?�+r
LHb�lt������=�?:v'���x|
�=�a{3�2��Y `X�h����X���#kQޟ��	ڇ��d'�-�Qx�@���V��6~>�i��x��c+�:�6!@y�tf��F&��G�p�V���80'K�(�1+x��s��?c�fDSH�[Ao�/������/m�����k�U���� �)�)�XP�c���=�u���9��:����}
?�>2Q��7�=I,Vu3N&����ňmh�n�v�v:l�i��+|�}�\�l*~�����w�.-W�"�q�Q���Ii�Ӫ����$v�)Ud��eċJ�:���sQ�̀������E���"���WZ���$��^�n�9E����6�dC����mg�@�p{�&�[ ���*{�T�e ���XnHp�r�#|)ΠِhR��_��W�aW�98��j���v�b�=nհH�jFހ��5NC,��F{�wh0���J���V�^���q�&������mag`��n(�O��=���BI���ǜ�8T�K�p��K;K�9�
.�ӈ�9�Y�I�X�&�l�oq�<P��X�w��&r'��~��Y�s|��4y�LZԤ�� p2���ʬ4J�u%/p�3���1�%B_�I�Φ�!�:�c�T���=]�53�3-z��ެE�J��ſ��˿�EZ p���,5������!`��E����~qZΨ���٠�z��W��tϣ�6�曐���Vssna��Q��E�C���?Q�LS�BḲzP7����<O�lA7�����i������Vx�[=����6�|�c��	��O�'� L�ޕA�Np+J
�l^4G�x,���!�8K:uez5]��mZY54���O>��$tW;5e3�~��1G�W��@��tCW���P���6��߄-o�i�&0����D-M�HF.�0�p�/~"�%ގ�����_�/"ܗ6r���&�Gh'[z��0���N��aCfc�1�q �[���y�>7<o�e\m�#TK��U���I s��������hc}&L~�K�Z�3Z$�iPrc��+C�0��g�`GAo�Է���)jbBkR�%��E%#�[��ulUUD�]r�eST2W�pK2$�i�s�J�r��pӖ�~?��FW��5k���^t�V������5���N��ў+]��X� �q@�7�GF���x-:�E�����u��w�M{z7��YgïUKǎ4�p�R�	A�	�����H3L�o��,�@���>}�����W�~\`�On�ұ�s�,�Kj�!�#ҋ��)d
3��m��в�����!��lۋpǰ��߽�������Aq��n4�,/ �����[[àg(5f���Ӷ��;P�2�a����x�1�����5@8�7�D`��ef�:8�/F�)#L�m)c�� ۯ��޺uF&@l���=�ˢ��r�ס���:]a��[�?nvH�wa�ߣ�IH�7'XEMj`ia�t�E�z�jc�g3���xY��7���F���k�eD��E�q���>?D��J��u)R�-��B����p<ck��<�Ѷl��K~J���u���&�<e�ZR���9��%��)B2eg��ً��!��.V��7��ϙh�dݏm��k���i����<���}@"�u��)����5s�+���ͬNr^r�A�0�w�?�~T�)�_�{m��[�� �nM��=;���ě�Y�#0�K�	CN~�����#�
��a���xU~���	{�m��@��/�|��*��ۅ���ܼ����u�Zn�5ҲT��Q�D��\����]!g`1e��C�L�����ݿ]�'��������*It9)�Jdg�� =���bdb9̴�	M���G~�!�g�T] ��nG������i��R��M�A�g��(�%���2���V�.F�{sy�d;����//�0��8'�t@�쳔�<���c���I��&|f�/�}�Wz"�Q��k�{�[�F��{����E����T��J���5Ǽ�I�_!9ARf]R�/�g=�>џX~$n&���+j�we���#����}`v� �3u��K��Z��q�H��>C;��1��ؚ�FA���\�o��̦ٕ�N�t=�gl7�8��ZS�����8/�0e�[��]z���}|ޥ�ܼ=�6Wr�Q���Y�!��l�>�	ŧ��W��+F���nh,MZ������.(�p ��h�]�Ƭ!�/qƾ�(QP����8��Py��.�H���蠖>���5��c{��S��e�)��n+�y��$�]���Cr(�{�>�Ұ�l���� �i�L�e��9s9襍�A�Z��XAލ|MѝW��r�-z�KDNb�>dڽK>67{�J$Z��Q�(6�$Q���o��4�eb��SH�~)��tH�Et6��2�-б��
�ꌍA!�Y�U��S;X�'��Ws|��kb}*��
�l��q���lk�a}����!�J��ܺ��	�.!8�;�^.�7�g~{�/j�H	7����s�%z����MG�=V�xR�7EU�́��&�^[�r�H��"Mk,�3#;~Mc��tIs�xVcz��&��/���D����S��V����[�	x�h���9��0
��J�{=�I}P����1�kZ3���j�����֕Ǌȥ����R��8A7<w՟Ԓt��G�Z.\�w�9Y���K��c��>U�9����=l����V���$��5?Tiq�FBi˒4�r��;,n W�H+��d�s���0򊐑��5A�tc$���0#h��a��;.uq=�Z��Љ�kt���U�	i'J��Pfӳ��$�W��^P��kI#I
���z�ͳ�Rv��*��o�`Du����<θ�-�#M��a��u6��,����},��.&��ʄiĹ��#���tcVc��RW)�Ww"�δ�cIn��e�\�8ҋ����	�G�nf�g��
��6��'q�Z���ܠ}f��A6(�ϔ���N���*l��-&*l`_9å!q��L���v�ca0.����%wA �v��܋�u	G �ARI���|�zہ������R�_�� ᆡ�J��2��*�{8˙[�X����V��	��bW��q�,p! 49R�:W=o�l�a�(�A� �#��2�Z��x.��N1F�?*1%��Z���H���R	..��	j�NۃC3��.*�F��1�Y`.�~X��w�ꗕ�Ec�b�Q����N>p<��w�ȸ!ǈ=Lx�a�Ao0q
jMrXA(��.;��e}ml������d��7���/�v�ҫp��hF��G�U ��c�3<h������0�_"���&)gI}���y7� .U�]�)�5����;+>?�ˋ��h�b���MċXy1�5�4���$#o����/5����u�
�EF0#¥a�#�A�Хm�����w���@�)T�py�8���#���pA@���~a�KN��ʞ���h*���W(p$���}��e�Ugt��`G���z� T��Pn�^�	v٥{��o-u/�%㝺=�����OY�j> �,��)�Gd&�/���f��q��ԔE1�/��v=-��ȃdo�+c�q5>�	i<K�L[X��c�UK#���)�娍�B%���c�tݖ�Ӭx��".�*��NǮ��G&+-��0��M�kk?	T���py�mvq�yѬ]zh��\�6��9e����"l�U���X}0B�
a��L@��F�9�Y��lDp�V1�5�r�峗_`Uo
bVV�6-�K�ҷ+�֨EwHp�)�@�Q?Bl#&�n�Lk�_,x�~�I��F>����!�\��Z[%u=H�h�q��%�NɑX2�uɠ%JH��V���f���l����,6��ȍ���])*/�G��G�g��G����N.�a9�0m��n��v�������?������HW*8.%kMNR�+�����Pdr��U��9��ِ_J(n�����g���&���[(ȸ,ψy�H�\T��z�t�9���`�
P닱C|3^���9ֻs�,>�4����K�`nӾ�蘳�g��C	��3߯Pt�e=k%+ī�=��U���H���a~\a]�H4q�-���cG�\���Di��4|fW��jy*���I��񙀽E�uFM�8?�ӱ8d?u�Ed��4����#Wt�w��c4@\���k�� %�	��ר��3�S.��~G�K^py�s"���/�@E�(v�B3>GD���@�p��� H�N��+L�J��&gB-���v����)I9ຊ؟#s��X��"�u'}jo!k����n�>A!Q��s��YYY'�x2���!����~}���"��|�LX��Ef��	c�n��������Skе/z���<
��Ѥ�4��/(���ћwc���;���D�b�(�:��G�*Wr��X�L�#����3��Z�R.��O)���]�9�5�c�mA��è���:8��������J������
V[]�Ja�=�X�̭[�Ȩ
��[�Z�ah��E�������aw#ޥӊv�>���^S�7��n3�Y"�B�U	����|�M��]��H��_\�L�G��1�� �{�����o۫���j���VJ͚�A
~ѷT��ZF��B�A8E�&3��/�Ͽ�����?���i�beX�w�.���	_q誅5�\�ޚh�e��nt�M�|o��\���Sa|fb3���q\@�ت|V�}õ��2�%�p"����B%�_	�.l�fA���.��<A�L�c�u�W\��4���-`��l�o
l�G9Y�5�`��Cm�<ް(�e��^�P&�S>ŵLq'T+J����f���#bN?��+6�ɗ-��M����	,+�%�k���C�$+D��X�'���g뉵�3d�8sp��<��=�=���^v�o��t?�^G�.��<~IT�Q߆*��e�
��Rd�l���Af�ju��X)���`���I7��*]G�/��g-\Ӱ���}h�`���%� K�<*��ѵc��%]��JFM�ǂ/�`\���N����͑���_{���/�`���R�y�wi?�8�P����������d]�h��еI�0��o�M+�8�'�y�1Vh@S�!���-�pn�gl�_=7���9��{��"~P
8q���;�����DA�s�� �O� D�Y��\�p�K�q�!I�<&�����9S�{�tC�4_�����qpC���.���t�D6����n��G�7�b�ii'ki����Z����&���N��q��i�)�B�h�h�hi�Ș_�`�<D5�r#�1�|5V*=�șP��b��x��>����}�ήTi�����d.���Mz��_��f�h�������X'�Pu�º��zIT ��C��I�ݡ�ڢY��`wMO���~gb�0;�>;��h��f�N�W�Xl�\���ݟ@��'a����W����T��>Q�ق�[^��� �Q'��xŉ�೵�(�~�}?(
	�'�iׯԣ�P]�>���MP��Z_��"�����~�]�w�rI7�3siK��\ȏx@xǒ���G���;�ԮQnIg^�M�jzb��Rf�{NA��}�ƻrsÚrTv����71�;������8k������G������1��Y��[�_���. ����$�k�Q�H�m+2�!_��|����+��oP��k��A?�O c$��"ٽ5Ad�nd�u���DY1	S�%�U�n^b$�����Ş��>�!�%[��������t�ou��U�>`��~�[�R%��j.
���f�ɡk�{'C�*�@՗� ��]��Z9���(�;�,K�T��}�1��~_�����]$	��ߦʥ�����ky�B��s�Ix��Ae��SEE�h���$v��y��4���:%�r�o�!�' \����R> �>��$�R� ��cS��T3u�.�v��\7ZfAH��3vҦ�}iz�v~��(�d�'ٍxy�A\�����HCC�v)jL�k����x� H˄ +
e�j蚗�����8<�B�k���M�u#�������>V>�K�A����C�ʞ�g��d`���Ky|s�JP��`+����:ֻ����V~�n�;��́jH�p�'l��*C����K�41����u�ܚ4��B���(�͈~���æ�D�9R���H(���V:j��?��������ӛ���:?�" �CKJBc���˥���-�|>�&V%��6fO�:� ��c���J��j���}ǟ�-�V �����1)i�Y�n�Pst,�8Q�Te��-������9`6�Vj��(-��bQ߀�����,��ݟ�5�hݥ�9�e�[θtcIX�#�C�H���ѡ���q��k�q���Wr{�X��0B��sv��7�\`����m,N��]���ƞ�1���:�3��ԳB�*����63_�.�$��37ƞ�U��]��E��:F�մVx���	��_��8FM�y� A(�m��!���u�8��8G��ݜ�,-r�������4 ��J�G�x���h�� c"��@PIH�b��\4�ށ�L��]bzs7=?�*���v!�.bU��10vs��|2�q�{��y�͝�,�%�װ v�:.B��b��&�"a��3Q�(����|oǁǉDv�7ڹ1��S��a�.C�y9BD��}��hn*﫥X\n6胿FlV(��/G�0�׍ZVtf���r����]��
����1	�X�b~`Q�bG�xD)/V��5��4���ҭ���\���K*����D`q�EdK_V�^G�p�����v�實���6�]ɼ����ᮘ��ğ/���(�❭i���8զG���ũ��o?����64/U|�s�8-eD���Ȣ��ׁ�4JI�R178��Ae2�p)��R�Q�������a�����Se�Vd�ߘQ�o��sL�vȓ�k�"�#�4r-p+�!���K��}�$%����Ckn ��p��$ �_#���Q���>c��-�C�;`���~L/�=ˍ�\)��ky�w�Jw��;�K��r����P!}y@�%=�(F���0W�!�_��/Zx�E]Ց�4��u!\.ۖ���qt=Y8͡Y�"�D���Ta�"w����ss�[$A���E�JR�L��ғ%�G�f�{�������#���� �w4�<QEO��TO-�zd[�~84���C��ڵ��'}�wV�-gɗ:��
�Ӆ��sω2�M�gF������,�p���$ex�z��-p� ׀/́�p
K��������K����X���J����:,S�0�A�j��Fږt�w���![sR+��`�}�t/�y#�2�|K庴���MK��[�����W��K�����F���2F��W�\ċ2�6cF�G؅���,&��
���+��fè�+!�08�W��,h�[B�K7v��l� i�����x) �V㞹� p l$lO��_��4�񭯃<��:�R��j�k!T�V��G�I_3���[���`6�c��R����'��v��'�S��)�P#����N�n��q�=��e0%E��⑪�+:E����O��I�"�J4<��٤���U�a��9�L&yMm0E�v��*�S��W:��?�_���
��)�رO![����a��.\���$r��S�Bn��P��hO[>y����+�q�h�JD�\�uO�?�񍗭/�g}R)�����@�%�_n@������~a� 4�M��͡ ZX��H`����� �8�
�$)�T�� �A"?V�mp����
-=���P��E���&��f�Q�E~�r�~@�Q�LXB}~xM(U�;h˵nGq)u���n��^��>���P�^I]Ek�VlK���e3ؘ�_/����7>�M4����QA7z���偵`U3�"��|qX>g�5uSL�'�dJ���[�.zAz���Rv�m� }��ㄆ�
qosD�V�I���Q��Y�4W�eA�m�<������8f�>��!/A�������O����ݴl��S:�o�)6��S�t��9�\[|��5T���s����ftZ�dy��0KOMt;Ȑ�B����T�5��H�p�?��e-�ţVp<h{+�����'.�L}%5���1+uI�	Q�vI��t�����?�U��طt���6�Y��Cd����!�,[�W\��/�S��qtI�������km2'�lasΥ�_љ�>2(���zX�&�
����Ҹ��ô�w��e�H��0]���[{'k���7����ۘ=�_	x�%֢r�����X256F
�*�l�gEc��V����7�9��:���U+C��w�>���H]Ud��E�Nx����t���N���mޑB��u�7���JX���R�_|��z܌���
з�91����t���-pU���S�d�nJ�lo�XL���,���kό�A����sp,!jx��;ă �38��Wwq/E�x����u�%s��J:�x��K�f�V����u7+9K� ޣ���|����Z�:�.]\�����0�jir��ʣ+�iL�r�4�L�c�E�v��j ��mT�Dy"����"��%6�������>�X �����9wXd��ÓȚt~wE�pc�s߉�i�
�tf�@GAh�:W����4����:���w����'qj���7W.3�ݩ$��|�^���
A)�о��d�יXSWx<�B�h�-�˕F��7���9����`���:`(����k��gO�1��D�~�� �x����D�������l�'��	�e��rܙָ� T�o�0��oh��2�MN?`��Q���}�UQ%���M�2m�,^��̟9n�Z�!c�F��_�ܨn�r˿��Yž2�R7��_�P�Z	���5Z<�yBԔ�x�V����%�!�Mi��5�{�wY���D�;{=��Sž%-ҵeo�4�<_b��*�m�S%͹I$����wea=t�|q;�<� úA"�΀� bV� S�|E�*O�~dI�a �o�\�����$<j�
P��g����1z����^��'�?0~	�h�`��S>���L�2�o�" ��?�с�O��i��I�<^�B��N��b���moV>&���� H�ǳ%q����SHN:��;ӡ٬��͌��ǼQ�}�i�ѵU�#+��PM�� ���78�9r�Nɼj��qJ0�����6�e�Gj�R��0�o�fJ}������yG�1r�=���P�}1o�jFf�dg�P���T?�t@��p�r@��f�~��r}wKy6���0C������%!Zo-'��ß���tD��&��E�)�g#!.:������a^�	�BYGh�ʁ�L�m����v[���!�g�c�%a����	�ګ�GĔ�>��܂�m�nfOP������=;�}�^�S����C���`�2t@�H)M��t�������x)f7�:�>J�W�oYrO�ՖǱ�S���~���w�ȿ�r��޴�����{r�)�.<_���ԩ�CΜLX���3�ܰ�:L�KG��6\���5���}��ݢ��?�a��&Ֆ��R�E�-F>5c�_���:����K���N>@�J�	���O���%?��֑m[�Gx�TI��O�[ؚ��z8��m�9pD������(�W�2��"���8a5C��ر]Z^e�,\eJ��Uϔ�l���(��Z�hk�o��d�dI�֩�7��0u<9�R:\zα��Io��������y��"Y���䭧0ѓ*
�r�@_D� 54Qs+��Y��s�#B�Ĩ��&jh�����prg�6UwZ(	���}��V�-���`���nV����J��g�#xj>N����Ǹ%V"�)�G�N|$��%��4=5��´�k�R˗��-{�H�d��L�g�Q��ו���Z&��(1%�,�=$��X��.�:�D�>��jy#�m~"����$��c} a�KG���1�x�#�btR�m��Q����a�/ٺ?�����.X�D!̣u�^}�X�k8�o���5�mK��!P�����p+�{���=�ޒ�N�(i�}L�]#F��M�:w�4�����wBa楘�gu��=���c�A���R�9	8�AAU_R0�$~���on��*�Y�̊��f�d]�B���K��S	Wty3Rq�(�>87��A�����y�� d "Wbc�O�ͪn!򦛴���,���
�ɚ��Nl�����2���BT�VSa�5x`/���5��ǫ��Zՙ����&F��C�A��t?8�
�%����v���`M��u�� �-�3��w�0�u�E�VСN'��z��ũӁ��i8H���g��/�8EL�|����|_O*�0 ���ۗ����4nY�0����>~���m��&meIt�E+���qW�A�ڠ+V�� 7\A����C�,p6eZ��;�xK�?����;(A3���7f�H�(��$�s�e⢎mc�	e����蠽������GE�*�a|�Y�Wi�7ָ�d0uh���.(�B �&^��dt�ݨ����>Ӛ���jp*G�Iqs4VOZ��O��i��^InA�>ΐv���>��9>]�l��~�yn���X7'Ʃ�m��O�w^���,�q�$�`���2��Y����v�&�	�6�Ch�4�-4���[~�:Xk������q'c�@��4e#Svȝ~�#�!���V =�1�[�uL��إ�7��m5+�f�㾑��,�A��R�5��T�B�-Ѹ�7���qSo ���z/q 2y4G֮�< ��/�b�OL:��Q[U�N.�j�-� ���dϓ��e�Cw/��ou�!P�p��t��w�/�vr+��2��|�]�˟�*�{n�`�� ���8�*k��<�����s�v�s~��ˈP$�"�erkf0 ��:�KW��$�pq�䙊w�g遟��+����e�DU�~ƃK�-TZ��˱�/\2�w5�X�b\�B�R�4��sY��1�Y^��Џ��A��|�|D�S���B��R�ZӀ���H�3*�?�i���!����ᦩ���L�>rW(8��j����E�0�F��c&2,���χt��1鈔�۝(�>�m\rMg��	a�y��H�Y�>@�V߾zl������	9;�;n՘70��n�g��,w�yk�B����B�n�)@{o(�G0OE�"���L���CvX6��N������/�{�D�u��^�FZ�.T��`(�}�-�#	�h�.�w�&le�pyc�Q��j@>����U�4�@THĂ;~��"��'l_�=Y�_�2�x�1�ͦY�[~L���Pba��.��0�Y�	~2,����wOc<���b�DӘ}�y��|Q
;$�3p�Z@,�PV�,{w�c(��
=?j��|��Bl���C����c���I�T-���b��?�-d';8�%�-��9w`��S���݌�ua��'P��,��h�6p��!����Q�:�nZ�r�k���Z��D���̅:'m�LO�f�jkQ��YO\ۻ]�xO"S�� n�M*�n⺏Je�k;_}�q��~�e�8����D0��1�8�T����� ��1Y��9� �=�'~�`q��]����!7W���rF��Qa�I�޲?4*��?F�
���r�< �cS��L��pΥO%�3d�Tk�{G���F�a��T���� P�=�jڢ�?��5%�[���Z�����_A0�q�Fd��0Z����"lb]�;��s-�I�;U�)f�E0fa<�N$�E�E�R{1��f��D�>����#u!-}"�V����	l��������|��P����>���u�ڗ�n�*\
�x4Mw���QϏ��$�,BV���P�c��p琦��e�o�klE�ҠC�Š��p+�|�t��D���5��m�J)ۗwWs8�?�>n���j*�Z]���3��H0�T� l�Q.I��@i��<�粜~�Q���{>-7ih������+	x���@m��GC�JVv�T� �~���=���z8!]�0g&4�v�%��P�VUb�/:���TՄĀ��a6�m�uy}'6�7s��+��S�`㨮G��A\�E��f�w���p��Q��N�@tO^����*[�� �>ћ��OW�[�&���{��^��l�hL�'���S$�z�2D������ɖ/�#ǐ��A{}|&���ŋ�q��)hs#�Meƫ$e{f� ��MDp�:�'��x���M �z	O�P�=<-�t�W�b.�pd�mA�Dm`���wo+/�s�a�Ŀ4o�����ڇ��͏�*����}�륥>f��l��o����9�RK3 �	r9��cSZ�.!n2���#��G_�Z�cxeH�uc}N��b����޲??��ۛ�\~�;O��x9���J;��?�,&�X��!���"��g�Rv
���U��旼,M��N�B��f���DI7z�Ʒa�C�1�+��H$.�������խ�ts�� 4Rzq)2ڢ��������}Zv�����1��;|+�*d��Cn����XW�R�2�ح�] ug+�@ �)��<��p���)��� ��tk�,T��n�&1���� ����G��4�z_䍵���1&�+�q��� o4�&c��N��3al�Rd�«�6j�`���vhR��BjPC��h��M� �r��c���ն��R�!	̈́�Ɣ~@�K�{8X�X��N%�M-ϕ����>U������B�G�C���7ތ��N���
�>�O&���s����ā���O<'�`ݪV��1VQ��hHir�PD9�0ݖcpy�wQr�K.'����D����{�,�۪�K�}o2W��vu�Y�#�!�x�./����������Q��&~-3¥2ӂ��= 3%�?7ٺt!�6��T���7�" �G6��Au:�˒��J�yF�}�:P?�K�����W+����W��q����)�ٿ�� �U_N��X��7�K~�i�BEUF�ʚ���
i�����[�ã[�hX}��q�:͇�A (�q�M�e� H�z��,�[�����c��dJ�O�	M%|�)�a�hl2��o�?��VJ*!�T)���@U��Ýeb�llF�+�Ī�#��p��9H�@,֐L�k����fp&��q��B-@r�0vO�fJ�w�v�,���=���жP#�uD���ɰ�(kW�m����kk��"nؔ]ML����h�țR0�ͯ��C)A�E�;N�4��6��ԉ��rp6}Ro�;[�z�,S��У�t�K�ϟ(��:���tu�xO���<��ܚ<p�[���
ıBf�^�F�uƫ�ÔMuHJRL���k��4? %K�cSH�ڀu��7�6D�s���x�#)���H)�e�>�ſ�{��u��|��S�o�m��5Խ��r�T��GY�@�0��o� e������c-W�K�@�®@\T �}�AN�T1~\��M���Q��J>�4�l�
V�t){��tm']����Xŷ|����P�N}�`�]%0gխ�JA�MZ ��f���s���!���z���1�iUJ����>�����:4�p~�����p���%0;k���Op���+��k���8�D���d���p�w.
���#4�GB%�)M�½���7:��q�24Ih��}��zSJ�u-D`uNpfp�*y2##�kzD ��U0Λ�"�A��P��W��R�|Y�p���43�@��^ƻ���/ͪ�8�h;Q�S"�@����������Kv�7dI�mh �Z�h�hk��o~�R���|�@��v]
	�s�lo����
�kP��&��T Q�g�c�bv1��H8�&���_&�ƶv�v�Oj�N�V�A:���p��:�<GF�~���N���Vf���:��٬�5Rb�	#h�I������Y08����d�#��%~_������Α���ާx�<��<f���#�)��AIJ�
�"���h��,����'��P4��d���횮�(u�_�i.(U ˬ�.쪄�&ӗ��9��g�������}�d�HZ��b�&aOb�����|y;�|�m��+ 	�l���?�S^>��^�F	Z��
�%�/;���Lη�]q
Ī���Wm���C9�!�5��Sv�^�ֶ�V���@������Ssmӣf[X"��m���tD�ݚO&-��Ԕ�a6�O�����fgF�-ŚT���o*>��!]/+WmTJ���w�D��x%�|�`x�H9��sͭ 5�����n`����ƣ^R�V�C�	��DV����ڷ �ݽ�I��KE��'���d6IA����o�����G5؏S�61ҭ����U(����]S�G)�C�p���a�g'C�+�����c[&1���k:wCez�D�\��?m�]�d$��{w�����%Q�YG����� �1��^��vꋉI��w D�����L��<GO��l���5��Ͽ�'X۲J1��V�bw� �O�
*�+&B�\v-�P���THhR��*g��$��<S�Prs`�%�I�����Z���3˝��ˉ���k�?A|���t�%����6�)X����
�o�������T�Ho��F
EZ.e�cy'^-f��kbL�Ӌ�9����IRt�Xqi7���P@$&Yz� �a1�J������,�}�V����!B��	�@�Y-�}�q���eFƾ�l`i(x�ʤ\�bkQu����:g����Kp�q&�/��ʑذX�G����<�Ƹ��YԊ2 ���������'l_Z��Qޭ�_�������B�N��R�,0<�jԓ=�9�9�0��mhJ���I�T��pN����/�nb��Ajp!yK�}�MX�K�]�(�j�4Sd��J�kT���N��f]f�Q��Z�L@J�
�����,�'�~Q�����N���/� Wz޴�@���Y��]�
v��
�13�/��1���`����2��o����)���hF�T�r|4ڂ߽����g3C�[|l o�{+�Be��g�ŕs8iN9�6�T�n�����Rb>�<��-5VX���)�R�{�;����H^zƱ�^.J�!���v�=�-b��)G��N;M��s�TLm�j��N[/�bJ1.��tb�%@�$�U��h��젱�sp�݌r��~1�$]$d9���dA�����x{V=q~����7��o��/Q����#��g�m}���:�	P��s��D�w��J�IBwHh���4�(M~�S��$vrK�H�ae9�x�@{<GiaMd�:�|�������r�>˿��Rdc���o�*�TG��b�� ��x��H��j�F�w\���ɒ.�y�,:<V��/��j��`�#��ٴ8gڎhJ��E�)}��J93���btp_�fLH�����/o�O3.R�㊧�}�K�gg�2d-o��3p�����j�	)n���7l��K0t�9��-��&/ܖ�j��)v�}M��g��zs>�t0��9-ؒs�z",���z�)n3���a���U4�3�����.{�9G�.~Q�>�Z��D��&#VP��G=���U�A<���2��,kA��Q��t�P�� ��lc9�ꋷ��=��	W�:~o;����2j%��Cn}��3���!.&:s��,����fS����|�-C�R�O�P�۽� Ҝ~D��g�����@�|�ݸ����)�Q���;#>1�v�>H��ً;3��A�?��d�]��d��D�kd�u�N��_�<¬���3c�B@�SO�r�jf�2�ь��M�N��	��2��)zy�9y�n�&���2�-�<����=i�&g�Y�U�	��P�����D1�C(H�/�;�i �A�aGfG�A�ww<-.�9$)Ip�<�2[4��{�g8�}ݞ��ڹI�!	$�j�_V�}Ƀ
W��jYo�>G�$47��l��M��ϥ!�:���$���Y�3�m�t�i�	���"vf����Q`>#�K�@��Jֆ� ~PK��w2��"@�u��xZ��5Bc���zG�S2���<�s
;���̎��F�Ϥ��c)�Ҝ��&L���
|{��⯇�P �s�����$��!��h$�
�6=�d6�d'�S��ԦU+���L���ؕ�͕صe���5u��l�O��Aa=j���(bӣ���u�I�D��͙��x~?�V���%�hEd��tH�Br���I$)9:�4[O�H`4�yr�Ճhl���,3��/���9ۢ�-�'�I�E�����F�gG�5@n1d!�Dp�[��\���s��R��o��(��UJu��40u��܀n���MӐ�7¡��3�cc��t=>�c��_�OE��Yk|��$V�/ȩ�( Z.}\F�(v՜�1�}4M� ��q����ZR�t�ea�{������D:,D�?'�p]��I����A�}��SI!-Bl�/ӧB�;u����o�u�)o�Y�L������7�i�(M�����*g�')/��50)��4�Z/T�fPh%y��!��������ܨ怗X�;1m:n�g1��7��Sfψ樓/)��c��˗W ���"��h�3�t�~v�NI��u~@߁!2��c�_~�!y/dNS�����v�Q��E�ɼ�qQ ��3z$Q�Q�	� ��yD�/3����"Ay��N���������Tt�ˤ)%IF�KE�|��s�z>]Z�k�l�����R�t��E�#�-��>�.2�3��=�)g.Kc��R=I(.G\����0�F���)����{F>)Phn�V�ѥ?`2���˥�gr�A�q�5!�1[��8N�f%�O=ٝ�[�{������4_�������!����EzI�pz(�>v�g�^�7�>���R�7�[8�1	��zf��5C�a�])g��l��
�>���A��t�q?��&9,G���N]�	*�����&S�X	G)���
��q)e�@t���v;��EԮX(ɡ�����\;U��&y6���m�N��Hd;��R�1�*�8��;�C���-;�3���cX�Fy��!B����8�D��\��岚L���8�;A\(#R��J��(�#�D���j�������zP�o��C��M]��Y���lK�	4� 3�>ݰ�y�i/x\��?����A��%U����`��ڈӅ?��y�j�d��!Ǥ����p��W$Om~��݆5�������;�< ��#���O�D٩eI�oJ�PY��c�9��4�U�ih�J^h��V�_�ԛ7=�wܒ[�ϊ��A�5�g�J�9yWϏ�WA}���q��0\^�3x�5dDO���kd����B��QxBq*yb��@C�b�x��l�0DY������R�_�����^��?~�gTZ�� �I��@eu�zβ���n��A �B�L[V�;����@������E:�X���F���c\y����W~�w`�$�l�nZ����`膣|��jaO7km��/8�#�,��@�d�ʨ��Ń[����u�@[0�ю�����jC�L����0'	��ҁ�����{z��f�Q��X�nI�(�#�	j"k��_���o_5V?�&�^O�!N���A3�
v���֞Ry���IQW���%!���%p~/C���Vڄ�8<Kj��z��æ�ɗ�s�ډVd+��HJ
& ۭ9jkI)@Ǩq�-�ψ�=�������*���h�Xё&W�(z�����%���H*:��-�{��R���)"w�?���g3.�[VJ�Հ��"�p�����X�c�b���?��d�;PXM9�۷���r�ƿXBe��v���7^�쿎kO�E��w�^�T�xE
&X7�����jE��|@�"���Xc��p� ���K��፺�2��$F3 ��J�l��)�u61]��e�Ɂ��Ω�QqVr�6T6W��^wփ��Z^�"E+@̧���0���/W�4���2�l�'w�k�=�)}D.+�Z�蕇���t��y^g��`���=ep�n��I;�O��ߣ�Y�t��������	��եs���[�FĿS�5�O�#�y���$�V'�Suci�3�����pg����[�PY-�le7j��4i�kIMj�U��g)�tn��?��u���f~�K�ZI�BI�N�OF,Cb$��B�Z�j9+��6~�[DQ���gՄOs2��BxҩSb�GS&	ssB��u���������-䶃���{1;�<\X������+�i�6{�i9dM�x!�����S�h�5�PbKc��=FG0n\�,��@S4B#a�{l��}����[�:u�T��ye'|�(y��/ɀ���9��J8q��CT"�ִ���t�dV4k%��f���:x-������>�HR[M�r+]�z�ANC�Kq�sx�8F6(2)�%	�7) ^���z T!{h�[.�4Қg� �ݖ?/s��#�Gi�$���C��O�c��2Ԥȇ&����Ʃ8�V�=^����*�k�P�� ˼��D1N+/{�,�AUX�:"z��?v�PR�a�
��E{yS���E��/zv��?=���f�'.�&-h�'X���q�dշ�l�}��"��ju�1��r�2�5(�Ng��Z�S'n	"\u�� 
Gk���[l�NoS/�.?1W&�^�cX:�Bz�x���M��Yǂ����.k����Q�Q�l�F�RNd��$��FY��ڰ(� {5*����)�(�6��c�;�Fl���Q�j����Z���Nybh�q1��W(��d4N�jaք0�x� �'�E�W��z�͐*�f6���Æ������(�
:Z�#Gw�^%+<X��c��������N�H|vP�(@���ag��1�=�v�=�W�l���y�B�$���jSR�����~��]s��;�ϖp��ӏ`�q�����c&��6��!���U
��]����R�a��ĥ(��/[�KT�o90���E�`�k�ݿ㉀��.n�q -���&g�=��{��ڿ�	��X�R�Ψ�C�����%ؿw��%�S����L'�]f�ݾ��cΚ�Ch?aBs��T�Np�~ur��+�9�A5y��G�������C����T??�����_'�y��nbq����c�)��'�<�R�o�2�n�vM�w�D�[~r���*ĳ0��_���+'d�z����/�͝�Y���8p�f����	r��KH�Z��4>�����X�����l���$g��Mя-%�i)U���d:�w����d`�c�[m�M� ���|�y�+�[���6��5I�D�T|ܘ����с"�P3Zj�u%.���+t�$)J@U����4��_[�}ũ�M�x�Aa�[��
:a�D�yai�@��o�]wv4U�χ���ŵ��������+!JB�?$�ѽ�٠W`�L��Iȑ�*��y?V�� rk�6Z�A �L�$����`�7�98-��Ĝz���&���fo¢����1b*P�i��C~9��1�w�/�,��NY�/E	�A߾>V�0FWR͚M4�x��5�N%��Qak�,[E�+&�0E��\ZI0l:��G�����9�١+���v��"ړ~ �����L>�N8عF�F�(�,��@����.H �gi��Ëế/�<H����6�!J��e.�#}��>f\�u�f������'6�A�*�aL��r(i��Z$,��v�(sZE��:�~zpx}9�hr6q�-�y��.*��[��AÍA��ɟR_���`��|�:l+��L)9(�jg�iڲ����w���,X�V��0l���i�*�7����+:	iȾbA���u��!ë����J��<�s�A��m7�����I�[gM��P-�D�,j��[���=�A�Lr"�a2���� �~�
u!K7l���*D�9�m�ΨM7?P�k�w��[���7`��^+���J����y��\&I�Y�ڒ�Y�����(#�;F����4</?�&lT5��*Xt���_O���e���5�v� ��A�4g"ƀˁ*a�9�/�N���dQW8�y5z����7H`��2N�u6Mɻ�-�lmݎ�g9�0�1���<�,�
X�/�>L�J|�8<�i$(�������)A͗z7t�A��hUO���
��{�am�=	���ݏ��
��z��Xv�g�2���}�m�:�Qk;�Vs�+�jٖ}t1�Yo�gi)F��R<gYV��|f0jM�0І��#�ܙ��.�t��z���)�=�^��dߞ�L�#c�
&#�U�Sn@�0�Q}�F�P�<9��?������7�� ��)"��!�-3�6@@�̨�3�����	�W�}���mFOε�P�����7h���
)��M�aKoh�H�ȊK�fH���c4Ȝ`֝F��w��w�,o��q��9���tJ��"�9���X��rڳ�^�?�d���~�|�͇}{���m$|��SA�ӽTj�ZنF6~<��x�jZ�C�Ǧ֝܋�w:@�T��.�\C�0M��AK�5y��~�,H���k�,OY<��-�b4�D�1�?iMԘwБ�C��9�hhLnjI���tNx�k�Y�Q�*���ޥ|�-�S��)a��V��ub��!.�������ae��L�dd3֣�l%Bd5t���l"�`l&�{�����Մ�������X��q)3�P��<����9�|B�M�s��	^s.Me�צƮ�<��B�aR7_?Go��`"��,�-I)���|�@��%IA�#T��#�oX�к�a������6��?�g$��[����`�;M�~ɿ�~8��8;< v�<&�pW�gAF�t�Z*�j���s��{k��&7c��	w���LR2V�ɓ�%��]ĥFt8�q�VX������<mS>>Yzɟ4{~*կ@�{X6�wrt`9?ڮP'-R'��?��$�/���m$i���?���,,�2|$$��(?��3���rnr�h:�c�E"�lٍj�j	��ul$���/��쥿����FT�l��d*Y~\8^6��)t������^�ŧs��2���In���v"P��0B������c�Ӗ���A�#�L���z��!�]��nG@�~&�s��Ө\ȭd�!�T_��T�D�1�&_��E�!��X&�3�3x���!�+~��?|��x:ڤ�� 0Z����,�gHulc�
MR��Q�2�h�7��o��2`)��ٞsl�)�����ߞo��U�j�;&q9R^YaT[F���~^-�yo���	�?����1j���X��g�Z�2I�^�SVAb
��mv�1çqS��<(���<��a���V�W��>���t�0_f_���tYX����qg���=����[Ɛ&8��녖�/?'�������~�R���n��� t����Ͻ�.���N�M���=8�s78��sP��WzϝU�'��h�{�������Z[��ю�U��)�]Ґ����@�_d��q�E��:A�����_B%��6$�AHŤ(��޷=�6�=�|.bc���,\���t{���H*R҃�
#��f�#�nR����-�#c�C�U�wp�]v��*��P�KTϝ�������Ϛ_���F��~�*�=��ǝ�/�"3=��=��P�F���{��	$H�����TS�E{�\�OroͱҖ�ﱶD�R�l����կ���q��Ap}�N��lɳϠ�=,�*�$atmy}�i$(X��gW8��~ݱ��I�V<�����~��FԳ���� cXyq�Q�i,A�)c�l@�ի��±�BK�a���;>-��돢 �Ϫ��|9rN/�[(��B��5`pވ[��������)�}�Hc�J��X�w���8���,�������2��/��(����b^Cb��l��8xoQU��X
p|<`�Ӂ�ə*�3��'�K���p���sZ(��DB�p��R�m��SX��>��\��,��7*�D�S�ٹ�L$����;�W��iQ&_�L={��<�VW���M1ۥ�A+x�9��{v8J�y̟�N�U��ݽ�(���m���Z�uAe�A���Z�W��w`�D1v�9����=F��@ށ2a�Z�{]�Q���Y������� �m�dS�	�$�ۨ���9��u����9�h̊�&m�v�@�*iM3z�r�
�P�����C�!��0Є+A����S�T$�ce}(竘�у����-:R�S�V�0Y�j�e��m�%@��5��vӖ(��<�/
��}S[��┖hIu�99���F��j���W6�T�G�2h�U{�Nin�W�k�0M֫f��S����VOL�AnH�/�SH/d�����KP�n���쏚�A�*��%v����.�3�;!����Q����h�^R�x���>Ῑ��t&7��sMM�dR4�Y��B[��؝t2�n�
͔ŉ��89������q�=���̈́=����L�� ���i�<N�m{�-��w�Z��\M���s�٥bazGk[�/t�)��-�|�NĽx7AF�Y�n��&��e5I�NΟNѝ!�u<��z�U̵;I��%���$�痲n�"b��I~f^��"��p�Ɗ&Y�c�`�9ti3T�Hx�����Y<v^��v�������� Ȍ=�d��ˁDj`��B�nFU-��v�%����,���5娷߅��e�*�2	ɰ@�"�(B���c��H)X����&����t�P*D��f�m�8�]����3���t��Щ��t��^N�z�i!���2��~�k�iǱ��p����/"��ULdKr�
Uj#�?6#�*���������aZ%��(�ef����l�rk0[��k���#9��U*�oQY�t�?��嫻� R��Y��� li��`���Q���"��{"�͒��K}��!�r�g2��$�Ա�T��l��ћx�NƼh>=�qG�0D!�٥o
�8�PHc~ڼ�.�4X4�88[H�!��W���z��@�l��	ɦ���ƽ���"��4*'�dQY>��k0]��6�o��U��=�k�ς3�83��X�(]t�!��^k}�p�kL��9��O��6Pl;�������R�*}8i�d���1;@-��1�̳1�6-m�+>g�L�Y>[�FLvC��&���)�%fOǇG�Kk�`4�WU���xc�C������)V?л/�����.r�N4�5� F3����C䵫(�����g��kJ��q��Ǖ0���(�I�u)��z,'K�w?����j�Fv�f��r�wB����}���h�ґ���JB��]C�Y�S�m���
�<��AΏ�Q�������{�J�ፈ%;V)���\���y&��v\�G�җ��aa��Śᲊ�� �;�fD�*�g���4�6W�W�.�]Q�L��}*�a���5��k[��$�U�L+��L��YD�]�AX�~������^�e�N-0��&�?�����SY����uB��"������юq�,[Dv�4�JϕE��+�������ܔ�W|��Z�kI`G�bI����ˆ��	i״�i��)�D<��0�=��=�(-Yte੫�D!\�)z����5�����<?~4�'��vr��mR��5��NV�h�<.`r�nz>	V�.ܤ�o|����ᰧ��Ɗ���(~� ���w!�J#�]4-
���3G�� 3���~�Нފ���5�X�<=�V�Ἂ�;m Ɍ61�������6�ԗbE�/c�D�6.�,_+OԾT��/�J�{e���s���)����6��̼.��sX�</�L��.X�r��x�Z�1Sq'\�u6-������v
ԛ��2���/��ɠ�JOM1��e|�ȱ�o�Iu���߂A�] d9/J�V�l_A�:*Q���/��΃��DY8c��S#rU�ݎ�+�VxI�߬���,3�%@c�ȴ�C�̗7���4�ː�����m>I/���y=Nͳ�}�K0:�����U
)���(\�VJf�:��'D`׋�J1]鹔�~+�b��r\w�{���Ӗ�vH��:P�u���ұU�����DI&,����fP9�g���b��ɒ:��Op�����$���V8φ}EH�A��������BvO;����7�$h`�!H3�~��g^lq��S����*Kdv�J��q���l��(�RɆ5��zQt�;����3�M�҇жT={�n25�n[����.�E�X�?T�x�d�ϴO�1����d��|KvY>�W������rC�Z���� ��k�Y�_��n��))� ������� 7~��8��vb�������������HC݋~dl!4�+FYc2�WS����ݡ �[��s�sd��vI��k�����l��H���⸣�� l�Ş\Ycj�n�h��:o�d��_�ݺ~���R�
u����&<֝���̾bjU�Y��=ސU��P2��*����j���vκ񉫏L����W{z5*r��W�6��:��"DZ[&Tg��r�9�"�ť��g�Try��`u�iW�|����"5/-�4�f���N ��n�zM��?Ø:2��}Yb�_堼�K(>:�� �h�݋�i�x���*ZVMws7E.K��迚F�A�;�|e�����
��>�g"�]��,w��^�_N�o����1�x&����L�5�%j��v�U�Yi�m�W���9��1$��`���J��\����wG̦��n`����]2͡�5N���o�G-������;r�S�Wڄp��]�J����G�5̕�I�-CXO��'7RL9��M����EweR%H��Z*��K[����v&B���K���V"�� �ѿ�����'6I����Is���@,��ڽ�n��O$ �ͮ}:�
�~fSF�h���Q������'��� �6t�
��KB�C0NpMJ)0XTv��]�@�݇BWvKVn�������"�����!a�R���W��	�$zȾA�zP�F}���:��)�����Q��O��A�����Йᵬ@��J���RY��P��/���^���2f's�˄��F�^'Q;��
c�b������B�*�?�R�/ `��� ��d�dI��sPx諙;[z4E�y�<:(�|����M[�VCꖐ��r#�3h� �%%k"LM�S����k� �q�Q�K�&����s��p�roι���	w�%I!7eٻ.j4�e�t�b���˄��t� = c�xCHI�f1�.Qe=��<�~���*|Y����5��oڔ�k��h����*��_�a�:�Ǵj�o��d�V�M��q$��.���������O���&5|�����J�zW������e>D�S&�k%�T�X۰y��W��`����{TL͔J�lh�m���1� �.|�H�+&4	��Ǆ�M9,mTb���Ġ��
��s�tj6�p�jX��nDGIF �>��3�	�����R
x;��n�*W�a�/�߼Z����է�6h�W��
 /���P!֖�3���z'�&	3ye�UPDP}vg���𢡊 [�Ux�,O7���]�-�y���pNNے2j÷2!b��@C�u��Υ2t����[`%c�v���hp2&\٭j;T���w	4z�.����Р�l�Xf��Ɓ�zG�:�T-}*n=�:�?�}���-���j'��v���M��T���+�N�����t�9�|���ވ+�M�6��� �F�m�Kh��桡�g�vm���~KsN>8)�8}����	�$;�m�� �3Ͱ�֤��6�א�.	�b)�W9v�r�4\�X$���_�������gkO��!eh62N&����5M˭��N}M 鑤=m-�6�Pm߬�í� q{�=� �+��N��7��'�Q|�%��J��4��JEN+y�q���|QA�۟D9L>�֒p&by�3?�`�Y���AԢ�tA7u�9�g���H�ڇ��>-ɽ�*�ڒ�۳+!�I}{��5` WH��w�
w���pG��w�rԹ��g	��&�`n�5�/�a�"B6u��g����p'~�p���®��t�8�)HE�!P�:	�sYB��S����w�Ђ�����a7N�\�6�|eP������o�%Y�Uwo��}y�S8A]�;��vలj����Ĭ
��k^�L&�9h��*7y&Z+���uJ2#e�Ӗ�vr.[��#��t����5�!�ƕo[,��؏1��r���c<�`8P�(u+F��Te�CC)J��Qў������y���n۔4��p�Y&=lt��p��r���i�0ૃ�'e�g�;G�Wtn�on�#���To�s|Lo�G�AhhbJ+թ8(��SD�w.����y~	V=����k��8��>���y8{�1r�'F9]�/��������@*
Cs���}|�Ь~'�+� ~x�(�´S& �#�4D���vl�K��}*�up�WvÔ#`(\��f϶�߱~E�U�@qԳ����c��?P�egO��b�lOb\;��4�ը h(Qeo�aS���A�&Va�C�D��>��]���w���Xz	cl��;/�L�9�va�`�|+|��L��f��J���8�G�r��&��.�9I�8�%�!��~7�o��<��_�ܒ����a���_�B#�+���4ޥ�];��m��S���qr.�x����J ���l�Ƿ���k+����sp|A�#��N�m|
	�����3A�{&\�e�4k���d�=4�2��Yh(�5	�P���ܭi��\d���tl ~m��{h���V
<��^���&��m4������?W�X<�qqd-^��@�x�
�f�T��$�%�H%��H�_D�����HXڍ�n�Jo%���V�Lg�����M��0�i���J�~����Xҝ�����nWQKϏ�q�	����}*0��im$����Х��jC&�""R0�I���Y��r�)�����n�@�����JN�Oz�(p���;�D~^!ZӺS���S��XD�<ע�̫���Q>�Y͟jq��]	t^[��a������$��l(�?��5�����T���b>BY�efP���=�;��k�i��K���8Wz��P�S��ee��p㻣RHH��/�q��V)͎�34�0�B��G�D��/ٗ�D��Ⰻ�9{3{z�~��&+�/=ά�� <좟8���'1צ1���1�o,G1�
�f
���'(U�{��,�;��λJf:m��?�뗏���cܸN0g���i6�D�
�R�>�؂O�Ko�3�<em�_G�m�g89�&�-���Na⸽������;#�N"�~I�К��Z�t�]�+���%���3�7˜� Ы�_�N ��*`��$�s�����͋&������ՙ����s������ʶpa�~BĆ����wY��F�]�i�*osu��v���T,ӱ[���D��Z����f�E^��\�[���x	�'J�g���$U&��7��z�7ʣ��$y�d����TVo��U�e����,�t�T��ьJ,�J��.��H�2��y�f��@!OE�65#X�n(c��Y%'m�2�^�X��m�]vi�G-j�瑯P�N�%�|��gֆ��V!�S8y �)`�M�7��bQ�?,��+�ڼ9&t?��y�����`A��.i$2�����P8��k��ؚ6l��L���/���ζT���� 8��^§�t�q�?�R�cE�\�����Hx��T���m�����E�])�~��fKp����>o��j�Q��^��x�Kb:���ei@cŏ�u�1���ԃ����3o23�l���$)'�PA��v)A��=�FM�߯7�/��A�f��c�S�}�����	-�Ҕ~��A��O����/Z;�lhEHb�|�Kr�b��Mhհ�a�ŧ/�q֋N�+8.�ܸ��X��t�h����H�VJ���c���#�đdͱ�~<�j�q[���f"�����j��!���bsk{x���
&��_$lw ���6�#)�]Yy<GJa]/ iw�/�ꅦ]���-u����q.󵐪���{eV�1��FZ�,�;�U���X�S,�󰾂�r�LAC�o���-��+ɯ����FR��ՠ�>��jP�mG��F+6��pL�y�K��'�,pfu����՛��!׍vQT�ա���H�p�R�E��ѿ�C�S��h;C}�u{�ä����p&4�z��o(X�Q��9y-��Ɉ�sY�l�C��ٱ�J�����n��-G���C�`��o8-o�t�d���0��H�k e�K������3B�;3��8��L����<���]�5�����#�N>��~q�aO�؎�Lb���6jR����-]�\Qf&r4s)/�������)ܷ�y"C7�XA5u�������/	�f������~��-Ci�R���4��(9wRjۉ��t���Hﾪ�����}�� �A'��"��|�~[��#����rn��!0)�m��(���*8����G]{�z�L�� ���{|�q�(�l$:���g��k�(7�!�S��I�b�m,���H��ur�Hj�PT����y҉5%���/�q}���I=�[0L_�ǭ[��Eټt�MEL@�胷�@�fv%̚ƿ_���A9 �HwW���ϖ~�z������������j�"�Yhms�Z�ib��� ES���I���ӓ�C�<17�� |9�{O�W_��g葬�#������c
?��̆�I��Ð��=���2��Wsd��z�M��AfU��?�p5�O��a��^��ŧs����4��9�iӗ��$s�{b�fe�	��	6��h��4��2������ K(���U�6ߥOm���)�a�-+��j�?wҺԌ�u��TV�(M��@�Zڐ��Q����d_��]
���Mт�oU���m����R�X��V�&�M�ʪ���E�ґ{�iUf�:yP�/�߅��~�L2P#�d֖��4C����Z!���C��Ť򙋿U*�$�LJ߁U�[O�T�J�7���Pٳ�P�(�����0��"f?��iGs��̴�`x�?�p�YR�]+��(iNj�Fe�^$o�J�B�7W~��֚a�|��e��K�ƫ�ce���5����V>rr��E*�i���P�wenN.rAA�Rdv{]��=>��\�i�����t��2�v['6��� �����xOƐکq3=��y��t�L�6������
S�i���f�<w�s�.�v�RU�*���~Cb���
�cC.0�Ǖ�P�5�d&%���v��G�aܥ��;��\ʜYQ����v�,@B� ���W]���S��!��w��rs��1��-�KW��ת���7�i�0�\|韁���ƚ$xz^�/q�7�)���<įF�B�t� �v��=z6E=.�n�*�1E�ϑ�y���[��e�ҼGΜ`����,� �/��jR�\�(��)6��e_Y�9Y�e\?#��>ԥ�n�3J��Nj��7-�tɆ���~J�bN@j�*�G"�&"De�&�3��!�8%{��ةc�l����٢����H�>����U��� Oz:��4ۧe����F.K�˵�f�s���^%�:�.�
g���~܋�>Z_����g�H�[�����SOX:���2ϋ�|�8�|�1�������O��N�v�8�}+�&i�j�� �m�ӝ�"EyyF��CbT�@�f�w�:f��J-�+a���O���,�^PāL��4���n�=ϕwn�+\W�G���s&t8ɒ�7k�h`h �b�/�|��fͤ��nmx�t7[Z�΀ϔ^{�w�;�K�X��/�)�?�/�6��Z-���Ve���]����Mΐm�_� �ޣ���{��V��d&�J�r:�+|�ƣ�}|�p�DI��|Cgi�l����^J���\'?��g�}��IT��������_x��$����^�f��줨tO0�ӓ�z�B����"�l=��vw1{~Z�<��=M�4��m���FÌ�q���3��O�u.ss�ش2^ik��1<拸��}��:6�)J�Q��*�A�c��Y_��8�<|�]�ӄ�~Lͥ�`�[�K�i#q�F�t��dIG�0��z�)#33	a�	�� |.�[/h<BE���?��$�"���p�ei�h���lm��3sS���,%I�S��X�D�zTWU��i�3W�e��q�ڇ^�~����c�c;��U
��69�m,>�~�c���(���WN�Q�w�7�������"K�7�_�Es3��`D5x�R��8Ǌ�&jp�r�P&I9�^?	r	B����m_��g�4-�r����eЫ���bU�x����0�>�z�A�zJ���jR�h��l5H��͹5z�ܑ`d������IB|s �	�盤���djl���u�~��������	����7镩�=aහ��p�ȟ�{.�;i�䉸�%A7�D|E���Yg����8�
&��3Y`��w֬WS�`8�P�YrL���zHg=3R0K-���E�c7Z���{aR�ڛ�[��r���u�7���C�Ys�{w�������!#̪�9_gt�.n3 y���o�|k"�n�\���ϖ��m��|)��}�3���b��y���J_O�6mv:'X������qe�i�[rC\��B�ȕ�"�s�����,�ĽX��f9��ci��r�E���]�<�zd�nv ��"��혀P"��i~'��8��3s��;0����Y2{i��U$υ�Q�t����*/�
d�Huw��k*��l?C�b1��z�������;]5��Y��8�Ť�p��ܰ����..m9g��V��a�[at��Ŧ�ә�]�[��/��L�W8���LP�M����2����S�T��T���z�S��z�"�06Y�m;)���
d��ֲ4h0�N��ɌY5U4qp�FZotG� �4�{J��hn�^�l%g8I*�rж�ݦb^/��sY���waN���
SvE��4��� 8�W�/��
����r7����p���y�gV�*QL�3�L!y즤=A���rl��jq��L�F-����ҿGSB4�Yp &�����Ƒ�����/ٖ�U@�ӱ��Y7�]i����INɟe_�?��-L׼R�Y�A[�@I�$`��o���LG�ԣ�a붿��.�}�
9u\=�ʾ��
	� 	&D^�Uq�!�(y��#V����ٱ���/	x;9iL��q���&�ɰ�������ɶ�����z��w�;��d�E�ڒ�_�"Ѷ�됎��R��b?ymґ�4���
�ȹ��{���J���q��®���^ gTHv2B�d��-s�@ƱY{'`��ó���T��UĤ�?o.g&%~mB��L�{`�.Ûs����sk'����������[LI�-庐�_�M�[Fo��	�E8.���n�Q�W��vJ���o���zմ^�Eٔ�{]Jzt�g���ta���V��2�!��w�\w���T�J��|2��8�Q�X��֗�mEч@M��?�Y17��D �T�g�S�K�El�W��䌊�j�JQ�e. X��K4�4lK�_h���7'� W����3���[B�A�3'�<a�'�dM���G�Y��)�+ЁD�o!4a�eӆK_e�S=~����U����E�]�]���p8���{%:D"�X����[;�T�T�F�QWe�ɜ.`�yXT,�:�����w��0Q���Q�㖜ؼ�t%l~�����~+ֽ��"�Ր�RX�	��s�a�KQ_��hu� �����΢�/�������ރy[),y]N���`Ů'��U��5��
R�!)x����WkcY��h����}5MLg�g�/��F���Y���VѬ�x�Nz����G��/�=K����u����#�B��2��jj�im�����,�Na>:[g�ʀ�b�Vd	(|��aܷZ� ��u�п����O����.90�ٞ�5�U����F��������$:�I���U�f����J�P�����=N[G|��#����I}��6�N�U�RY9'���M������
kگi�4��a���p�(r��|�H���7d�C�N<�)mq܋���_�����/���Oj���VW�]jD6c-�E!���e��5R=�!�Y�Aі�lؕ�G�]7�ԍ�jR-+s� j�H~橱˗)3�P�#*��8t�	�"�=Yo;? 'ٗ+���*�K;p��<��/�{:U��>}���q_>���oHbP�a���yc��:d�"��÷2	F� V�-��pqZ/�Q�Mk�ձ��ۯڢX5�[�G1���g�[q~�;��؆�3
_Z��������BF���;�8�b�L���-EtV`
�*��L6*Uf̭�p��!1���d��g��f���&�B�̢�&2q��r��i�D�� ������_�?��%�d��DXw���C3a+9����2pN���A;dJ�.e�K�EToyWs_������q��Sʞ�R#����RЦ1��B#U����ĉz��u��0��j޶#�7#��w+CT��&�#iܧ�
ʎ��:F��v�ؽ ����D�fqv+N�|��L"9�3��]͊��x*���݈!pd�"�|�/�Z���gm��p�NK�v?��f�Bn������)�e��`Y}7�k�on��"}��J��u��,W4���A�o�{S6�4��ӯXFMy�V�Κ�󗚷�2�X�ȹ���Ԏ��&ne&QX��ˬ��Rzd�)0�9��z�ɉe0s65k@�n������V+ޢ�6�{o�ܖ�N�K���]��f� �]����&�7pN�qB�؝�x��J��^~�S���+�[�
z��x�DwZ���`Zt^�E �9YAE�7�e���Ok�X���"���?k�����Ʒ��� �~�� Jm%��<�Ly�0  ��g�x�=E�.L�p_�~�����q��u�"&���q�୶9B.)����@�ZnŠ8zg�&!�Hݴ��]p�?�qp�"} ��q�e�H.��"pn�a�������;�{�cm:�>��a!f,��1�⍦��75m��_^b���c �)��d|̒�z���L�72o�4 չ:c����#{��Ӯ���W����;� x�6�v��q�WB�q�A�!a�����0�e*����M��Xƕ�rCs����#�΂��a�����|�]-�7_���f���D�qғQJ[�t�˫8O���w��Vcް������}���.>n$�Ɇ�*!��j�Y�~Mo\ ����s���UV�2���i�����/���}��^m�B-2������Q"���u]Z�S��)��At�y���\��As��'6�}�h�:l�� ��I�gd��I�~�8;�Ұ�Ǻr@�ф�f�`@�|�N܈����䉕�8~��0�`e5đ��b1(��q��.��uVja���fހ�76I.���c�6}�:r�� n���Qs_�xqAc�Z6z�ڜk0�IJ�+�~�+e�wԐ�$&�-��a�P�=sXH�l�Y��{��$
�C
�4CNo?���"ܻ	�����`N�2��uD�h,����]� DZE���������n��c�2�B�W�#(�B�Y�f��s�U�#�Z@.�թ.�q�]*�4`��H1Js��wv��J�-|��yw�+�s!�+�!�Z(NkAX4��gg�0f���3r��)�[DWE�}J�´�;���%�yp<�԰��S{�_�9Ţ�)�{��5�"	F0[î�:�} ��"����4U��C}�^'�:�m�[�2u★�Ի���h:�T���KZ�Wa?���Z�)�����p	l��7���#��0�-l���r�$��s0
 9l�0k����c� ���á0�$�-!�+�N���@�z���hO��X�w��盅����W�^�

������.���i�Y�$��_�3,���[e��4={~������6ȯi���A�������#{�X&�+g�Y�,TL�+�+3o�m�'TT!:-���ͣ��@��Ӊ˾�ٞ��_�z�Ү�bx%�`5�J�w�y�J"�=�]���� ��=j,$�"��2�ʡ��~g�Wc�A�����Ιkc.L_y_�d���x>?-g�,�߷�'����s�WB寛�֢U� �8�V@_L�������< �E:h~n�WD��n���?�q=��ug���_����gѿ!qc��#�8q��:&#C%b8��dl#��;�zG��p��������9X_������/���s�Za�zU�T�K��L��L.��9��9�u�Um!�'�y'�u�HGM��r�a��	ۖ���H��s�A�a���(�'��l�Hk�Ǒ��In�uk�F*���JLSCӈ��̨{�I5�s*��L�g3����@M��m����O'/ J7��������b}��;bJ�FMD�A2��{���y�箙+�Lt0�A$��]֚��d�5͞C����ܤh#�m�yw�R�d�؍+��D>e�@utu�/���%����`���7H��:����)����+�aغs��~ڐ�����EF��$�Q��^4���h+Gcy����T��0q�t�e�p�WW�%��U[�C8�&�>��4�5��Ŀ�����8T ��J�֜�U����kή��?��y��QXd�Qi���m{E+>�1~���i>!��z�>SGD��~�G }畟�zdx�K	% >'t�=#����˚H����z1z�ޚBg!��傻�I�Ϻ����|�c���}��UPbh�����[��T�k8|�s\:��QkII[�p�]���0���	?��Y�ߧF�;'j�}�:�w���#vRoz.��^|�K3x����jz�x�·.t�)M7a�7;N��VϷ����-�v��Z��X4z��ƴW��m?��`����2kӋ��n�󚓸 �X�
2��}�X��L�`	�,T��(r���:�+ʭ^���Nį;���=S��E\�Bm���PU�	��3��U�("��Ah��\),|l��*
�Po+/��R��xU��G$��]�a_����T����a�
u�(��m=���L,�aM�����P���oyK�E[[�-u9�Q���\"/��nf9��d�Pw��<Vj�sI������SȨd��!{6 ��_ټ�G�_��@?wo���@lP!�zG2�Ut�+���'ΊS��8h��q��3�NNKa/}� �����6��K�*?7�vK|�<r9L�8��mM	�&�L���{�-B_�xB�Q���|,Oٺ<������9��h	���t�#���-u'�Ը��c�A�Y*��E6T!��MZ��d�7)��^�&;�To[�����~uH�k���F��q��q�&��
�@�����8Ĳ���m�߫��f��՞�O������3׶7��II�(
�u����E��C��iX�����X�-2~�/�Fr)��7sBT��X��+�(��f��C�<�/����]f�n�N�C
TNW�� �f���7��]�1@����J�G�?I��l�/fU�gK��T���G_{�c���o�oxBګr��I�~Ԏ멻���Ϟ��[q�M��V"�>Y�^S�F G���A��G3���#���
�I�G#����F,�ɓ��Č<�^r�k,�oF���T��y�WL�ߖ*���12<��U�X)EZO�������M���`�ތ&��Y;o�%�e�xf<u��0I����I��}r��Fv���&���I���q��(��(h��� 
\�5������7���`��(� b�KA���2i@7q�dM���`���*�$5X���"��ZJTr��1"�[�N�{�;�:��U���B� Đ���������2re[׮��qL�;\S3T*��u�˪���d�l+��x�������r*�o�S��cz��8>�',)p�:U2��L*)���C�z�I�͊��%�u�S*����/\0�V�����p$
��l�����	ӓ󆎕J�P|$=(%u�p4h��) ��KT��'࿦�U�s�t�r�P�@7��M�c_��-A��S2��9U`�O�zՂ���Wt�5���y�Hj���[��.OS�E҃$-Y�,JA���,�����XM׋��APId��:3���	�j�P����ǅVU�[Mg9�j�+����l��J��R�!:�_V[91Cns	�3ԡ��hwO��q�%@�;~�e>��ǉ��{�\�,8o�*�^�tjδw�����6`V�*�K���v��Tl�ٳ/��|-���i�as"�X�O�n�CaF�����o��7�#��{�q]��T�DQ��W2n�WT�w���etIgqŹ���x������³3�ż��s�h|�ll�]�.�&��i\��%F�]�Aѓ�����\��o(鹹����T����/
����v��##�Q��E���Qh�a㕘Gaկ@s��ϳ4�
CZ��i�=�f&�<�hy���F���F�j���f+�	��[xL�zX��[y\�&�纓�M�o��隵- 5�LO~t)��Jw�̖s�k>�u\(λA�mw��C9+`s�c��錖��"���`�
o~7k΄Є5��@���O��s���sP�E��z�*�_�FQ~&�p�ў����S���Қ�A3B���FZ�cU=����E��E[������ BÑ(����\�swBwV�V��3�/����J?�ʡ��4?��9J^fE��w�c�[�z��%��p��{��N�Lfv��M���Z�ʀWp��o��閕��B�D�0��QtZ�H���Y@]��>WT�����0��,��d�4���w^��z�0�>���V��tni���,���>������2IOkc����b�.�P"�����;����m��Z5�z�v��,���	���%t�V��&��f:�lE��x��^�>��uw��7���G7ht	�����K����Y4��JM:1O���X�ϣ]���*�Ȝ��}�y�"f���D2�h̆�&�o���eK'L���?�iм�$��x��l{u��~���>wضv�{��N�q&0u�	3c���ξ�>������95C������!�4>G��q�!؍�
��)�{@�;�Q�0�K��Й?���ض����o�a;�c�2ޥ1�C�h���M,B<r��ʖ��ċ�76B��}�q5�k�:��@�ە�����0<�D�����ڱ�r9���\j� B��vN\	R��sF���u��`Llz4�?W�e �˺?�[���mYMl�A��� G�D��1���;����S�R-���yո�������:�֝h3,�š�ݗ����1 ���wq�\AtT@D�QYH�C|q�J�ֶtk�0Ҋ`+�[N�Y�,7-�Q���x��4�S�nR����
������c�Ch����^*&Qr�Y�)@7��*����Y�_��!��l��r���e�UlU�OOW�<�nl�{^�ge .��=�lS��Ys�o��Z�b�xؗ�ߌY 8��_=���k
��hl	�D�v�cy��H<���\����T�k̮Y_ن��g��TQ��?+E�+(6?�����^�Q�`��KY����~���|����v���7��5���A�kPEY��Z����&�e�dE�ёᙿK���h����:{�q�V��9Q)v�+��9/��mΨ�Yݓm��^x�wE���	k��lϞm�O�ؼ}!�҆�"�T�� ���[p5)����8�X0m4uz�FE��y����r���+�Y�2�F9� FƧ���xgCT5�\P�Z�$iZ��3?��-�I�Yc�u�
*n��e�C%�6N������Yi4(}G������`��:�J�J�kl�;�ɄnO)B�Ua��덠��nc#
-�i`�V���9^��}J�&����MM�q����Ss���G{3���>N!�HEQ6�Ipm���}:�"RDm����c:��/u`��B"yERP��B3��F�
��dJE	Q԰X���2a��M�OE	2�@���n��- ��3�<	`ɴ2,��}bLF���k���"H�P4�e��Ϲ�C��B��L�_�$2�SS����9��-��R��¥��-�#��m3i�O�#��$g��-6�q^_1Ȫ�c=cf�^9V�$�	⁫�ֳZ���AB���rD��x؜3��1��ըw�&}���6J�K�o0F��CJ���)��}Gx:�B�o�!:�GFی�k�D������dJ	hM��L����F`��Yg9��L�*$օ�8����������}���ÑBB���*�_bi_WO�LC��~W���hif�#�|x���p>�q����V��?>�@�����?F�"U�ɟ�B��03�5���T>x�5��`�=���E ����^���o���D�,������xڬ&c������r���������n=�s}������)�����h������p��~��wUa�@ӓ!@�F��95��Fcb�^���,6�L�[D�V���q�Gf��x���z3kHv�z�	��=�l��Բٖ*�y�?�S�|��PQR �7MrjX�:G �L�y�\t{L`)��jT�$�f��ط����������q��_�D!�s=JR�i�7�1d���PR��k�0S��Q�'��&��mj�%:����*�Z�s��ì��V���sO���e����5�!n��7@Q��}��I�IϩgԦ$���ZN�!D�.P���#	����8�S>�T��RA��1(z�<�9����A�,?R�G�G j["<-�oƨ0�^Ag6�@��6��ɡ�,$�y�_Ԙ������0�E�lZT)�y0��3	:<j��7��6�o�(@m�&k�Ct�S�1��psY�j�{m_���\�7b$��ڡ��WY��i�]]?�� ���X��E�� ]|�>A�_y"������:A�dCo`E,Z�TM�`��w.=l�؛@��<����)2�?�ؒ��²a7��4Ft$�>[�ܬ[�9	[�݂<N� *��ex���8��Q��Z�?��W[����TfN磟\�ér��ھR�$n�5n&\l�ꆫS;d���4H��k\���}���е����l:=���N�8��'�±�l��y�4Ӊe����9�rT��t[R���NT���/�k�7ӲŴث��Dçg�hN8G����۱��M�]U�Vj�!���x�^��e�"�T�)Ɠ��;*�n����Ք�EmV=�����C�1��0\�w�j��'��P�!�[MH�J�5��ܖ  ��T9������5��#"�Ԁ6L�(� �ZUh�E�0��oR�u�z�c�A�J�oe�-#������t�$��3�ܕ������������n�h>m��e�������`�ʣ��r�.)���L�D�G���H�������{��bӳ�Z���$��Z��B# ��@��	�-,�R�{8-T	������5̾\5�ߵ�)]{}OD���V`A�׊y�ϯ!U�ac	數F��Ͼξ�TI}�2? �_�iG�ww,
Z�RJ՜haU���@�(Ϭ���s�jߔG�Ӟ�����<&�s�b�� ��	��������̷&[�ĝR��q�j�rN��i���;�&�p�)�n�Эڡ�J:[{�[P	^6�+��j�����YDP�CHn~�,�=t�j��$d~G;�V����k��ť��U���ج�ob ҆�zҟ΍t/�4�FXf������^�sp��zB��'�rJ�FF�ƍ	F��V�~��f�\��jۈ<86ӝZ\]"�c_��_� Qcc"%����
����[��P����y�1s�������/� ����Te�R�/w�칻��R?�\����y�zv���h	���U�}+������.q�!)T�耜;gӚd](�B�(qE_�<E�m��{V/E\ګY>��%����"����l�?P�d5�j�ێ�;M�wa��0�֞�|�V3R��\���B��m��Q��XZ�Ku�lr�97���vm��F��]��ܼ��  g���t���ϫ0Gʋ��;�x��e��
ޖر���[��E��b�P:_�miM�R�s�mo��D3��Ć�H_v@p�<W ��pc�yw�0p+/ı�!�!�<X�F��<ö���E0��K����¤ۮ��C��l���Z^$��w�'p�7�f����I�F2���h��Z�5�EX�i��	�o&�+�(��F�N���H{Qd(�����L�z�UI�:o'"ani��h	��9����[�x�����d%�m7w�I�f����"Rܜ�U3'�9��3�D�e�#칊L��6�Q�����+��)�Y��hH� ��$��H�A����qO!�`�k<Ov;n9�%��tk�b�O4'"���Ij`M���;�YSw�5�RW�' ٔC��� z?J��C��{����G�Դj�{.+cH���]bQ�
�1�������L�[ş�P"2�)�4G{�ԥ����fy~����\ d�N$�P�t�sw-GO�@'Q���Iќ���a�uPRz�B��=��O�`v�B��!U%��T��o�GYV���Uj5��eeEH�����z����d�,���އd<ZW�Α�E!'�q��DhN| ��1��Kr�o�F��}��R��?{_���E��m{��>��t=#�B��G�fQ�>_*5�����Q�p6�~�t`��Qu��fM�?On�gzЉU�jB���ź(�إ>���rdM?�3����)�Q����)U����A��i��ڙ�Θ^	E��=�����^�3�3�p	>��pWf6K�a����X���7)y��Dj�B'5d�D��/\��o��sYE�q��U4�|xNą��3r�]I���"�
� ��:&�F��̯��'S:Z9>h<ٚD�`[g����_,���\נ���	t]��d��[�2[��V�ʇ����N��)��1��ewi���Z��ߕ�܀]�-hnm�N���q��Q��T�۫QA�8�%�ԇb�m����LY�ߑk}�%���>���¤�K���s��S)?8�G%!�t��
re�b�#�.�*�C|$�E
���
��;B��	w��(�pfy����ݷ^��Zv�s. ::yx<�r5��q��)��2�A=�{5qn�ᜏ��'N�8\�A��
������1��Z�E �����9����r��J��jz�dI[�"��E����~n��ы��R��b�:�Q�A;�b�5�!]p��r�)&8��9�ة��jɡ�F�����J�y�N���v];��A�����HɛrF;��C���~�񴩏�;��>Mf>�"�������e�zuԂǠ�g�r�?�_~��2�S"/�(;k
t�"T
�31I����+���g��_�t�J���9�bGYO��_��ڶK.uumQ����ѽ�sGgy'C/e������A->�D�힌l/6��^��"�|���Y\�h�@����g:���@?L��q��$�`�2���k4��ď=�_ot@ŋ��~�J�!u}։��K���+C�w���q;�t�,��{۲

7]j,����aI&����Jl3���	�3�$��������ᣌ��)M��"z�ހD_=�ְ��62����d'���,N�}08��<�פO	U]U3�wŪNmn��g��s�X�hz�45������=p��P��;�X<�$�HO{%8'���}�}�wT��v�E0eҺ1�83�X�H��8��a�9w���ŉ>�w5^�;�%&���7�����3�8sx��Ф2�hAp�"@�p���\8:��?)���m��)�|1E[
���,���+�cbO����s�~5:�xq��^���)Y$�-Va抉��꺮�e��?�n#���y���a%��_3Q,4R���ǄHt��U"�kqf�̉���= �$�Wa}�I�C����~�@�]�{��C5��pď.���5Ȅ���OA��.a�(�J�J��-���}�2j���w�vD���<H�}��N, ��BGG�r�Ĭf�!�Mc�K^{�?�����ȿ}������P�F`ٌ�$�$`�Muz��%����A]��o����U�RIm�Z�d��Nn�õSC���2_���@sF����@���"�2��ڈ��	��Q���F��E������s�#y�jw�]6[Ͻ�$�qD���	�+<��qu�G*�/��Gnp���Ȍ۩���W�t��W�W��Ery2�G�GA_�ľs����*<�(�I�l­_�H�N���d�;���^m�"�M��~I�D+u�M�}���!�H�:�]��͛�$���sʿ��6ohw�tZ���� ��WE�0~x^��j��rv�x�t�/�DٍU�E�K����[X�w�f���%�H�w��P#(���/�k��_RWۃa�;�״�:�I�-"���	�#�"�h>�\Z0��m�#2X�v��b�겭���P^��M�d
�64%lmRT�Γ1 ��ʲ�7�륅&���%i���a� ��py��:ܡܷ}����]���E�{I�8�XNަ�t�q4\6uP�f����0��`���N9R��J`��]�dr��>U7�)0q�=�٧�Mv�M�vXOq~I�z��_D��*�c$ǹ�ژQ
�³�k��8���ۡw��3�>�y{h�B	Hz��h�q�\�r�]�/�SO��j�֡�<�Я�^h�SC���Lhw�	hNz�Y[��r��=���D�.Y�;C��s��Y�^Q �a?=J�.�S�/��jT���K����2�[�Z'��A���J���+����ֻ��,�&�����vi���4�B���2	՚��/	�B�
������ﻉD]U[�K`�f��������Ύ��Ff��:^����=<V�u�"�퓁�{��}e?*x�U�r?*�l��_[���==������IVk�w;��{�(r�3�6�žD� �t`������	R?.!?�;˔t��ϸ6�#!�ї���Y'Mq)�q��*	�g�a�'�< �Ŀ?Q����\�d,���(���%��'�.qΊZRu�q$��{�-��d*�g?�S��v�* ����L�ei#X �B�%}Gtw���Q?���ph�30��[A�s/�j��0��ճ� �~�8q�S���P�xq�j��P���� ��F�./�P/��R���=)�8��.U:Ǫr��������:I��X6ĕǢE	�X��#���ւ�"�LUak��
�C���+ ]j�g���Aq���(!��b9 s��-+D��>LB,2�v�C.�T�-����"˵\�t\,�3�"��8��^ܬhSЭcr ��a����n{�)8�ocvcZ�qk�G�X�������lbVkV͢���w�����r�����N}��2��5�i��'�Tͱ�J�|ZG�FNKp�z��,��}=|:Y�fU�]�a�n���:鷈J;�CgV�,4���҉(�p�; юx��ݭ	��L�,����Ef\�d����E��ê�s}Or+��'}��}��ݳ"�a�0�e%��VA�}��d�Vӛ~T������x\�j+0)��� Z1n�m8����K�^�Ц<2�"-��#���3��|�,��`?ś�VV�g���W�Te��A�i!��3�i�ڙV�[A3i�K��f�hd���tTO��2��;A<E��Y�~ 㠒OǁG�#�Vahce`}��6����E�
H➗��;:~#��Mc�GT�=j@�ٹ�Af�Rq��}�O�|�a�����dQi�FT�����C��k��&�3��x)6��d��{����"�>�4�
9�L�5�����Q!�{�V���hd-�o$!����Y� ��|w���"3f�5�WN�y��n_M�LZ��")�� �*= v�b��1��~-��LCL�Ȩ��]�䄨6&��/�3(��v6}Q�������t!s%!zB��Z��D�>l� �~�m!��8��e���l�ҵj_���~�O�\&��Վ�Y=�Q",u����h��t3�J�!|0�2�x�e���&�$��pr�(Vp�q� /N8D�\8�\�gi�#+@�	Fr(�<�_�LQ41�"A$��mn1�!��\��O�M.?{���\�����8V�6͚�;�b�v��)
~�z|�崖�ĺ�� ��p��3uO.s�R�_�;:X��
�����e�/R�����e�U�?�|E���H>Ն)��[T
>;�C�Dϰo��9��|������n6if�oM#g4�g�}�4IS-�b�s.�E�r�3��Vom�6X�p�����Pb�
7Xz������T�@��E19]��Lir�u�c�m���D���Ez}f~"Ts�r���e����&�����)O�SG$:�NH�L�x�n-x��$W#��3F_ײ�����_	�������|X�g�;�  ��{�O ��|7A��ć*4E]�_0)ʤ~�/�º<���M-���呈k�AY�j���W��ղ�t
׸ h^�^r�-X�u����[w߷��*��4G����T1_0�Ġ��v�����Т7*��P��I��?I7�k�^=���w{义ǚ�p�:3A��G����?ϷkѬǴ�qA�x#ɯ�@��F�O�C�4V�H�+�F'�! ��7�X�� <n�[�q(�ĩ/Nm�8�Qb���v3NI/�O�F�7D.Җ�f���X�����\�jh���ӧ!��_0_X��2�bd���{ti�/ޥ�$��Dt���e}��@�%G���
�����t>��������;�C,�s��=s?:g�;�	 �w�.}�6���>�$���aڕX�:��E�[	¤�!r����sj���j��[�� ����Y�V��'�y��ޮ�V5%xJG\M\/�]�ŉZ�Zs��2L����M"��O呅;_����h����h/�H�@�4`尴�b���я���s���p����1PƷ��6f�V�+,m��$�S�Y<�±7*��ŧ�%}�HWX����9Rt`P��؁Zh��?�')Bl-,X�ּ��^��>��5e��Ћ�OKhy�0h���d8��%�]�2�0H�z%*  F��tiB��y3��o��ު�~�|y'���{d2���ٯ)@�S{pj��@O�c�X���ɓ�I�ʁ��� �X��V��|�wp
��y�!�!���-�Lc��4s�x-}AO�6���]/��ҲEn��K�*'�7�q��w�9������[�t�& ����6�p�2��RM�
�v�����^��- B�WH� ,���(P��G�'��*HFʼ�AvA�2��%r�;�x��D�"8JA��3����-�����.AV�.h��ӿ�-;�c�����Mí������jl���*��>N�rn��~0�D�)!wͼUf>Wۉ�»�ʙ���%7�B?�8c�1��ݍ�N��ay�ݞ�I����1-����:{�!㑨��GQ�tw�i��p�\*1�+A)di5Q�O���~�S�l�D�%�%l5'�&�'�?Q�N��*�Ta�;K�P��w�KH�=��&;]�;0Y��(�D^�?�4l�˜�j��HS)�ͥnC�m죴!�ح���#��oM���b�?��/i���Ėxu\vl޷����@����y=��}��?8��ħ�4��D���A��?L9��ȵ�hP�_Zd��)����x9	�eq�hp���ئ\����j��_�_�:M_�F�;�Ր��lv����� �����qrq��sY%d���R���َ�'�%s[�/�Z�ݷ.��K��<Z�xX�o/0TP6㯆�Dՠ��ܤ.�Q?	a�O������:3�v��u~K�ι������Ǯ��G�6��YȻ���d��L���<����S�a��]7S�y.#J��qt"�h������㠕²~dA
���>�b��9�P�m�8��v�I�eڒ3��on����2�^�b{���0�F�[��������(U��/��
v9jͅo[}Q�k�$�~���~؝5 <�>�L��(��1d�8Rl{�]��8g.�@
�_�֣�i��\;�yB��A�k�1P��|��צ@l��s��/��~�pn+�2ģO�k��q�K�K=�]{�k�=lΛ��'7�[�2:B�/3u's�g~�:�!bR'l�(�`@�F2�jѬ#��	n�P������I	8�dTQ}I��V�����G�R0�T̔�#�"8f@l�%��m�[�B�>+�[����0���n�D�r���� �W~��״GZV� �lkmQ�B]��lj��{�-`C����^��V��g�cA�'���w��G��^bi\�cn��4��g`Ge�a<
Q���M��im��I:��8�h�����^<bq�Є��� r0t���v9f�ܬri��(_��� ���Wd�X�"��9u�1R�f���a�X�?N���x��&w���Ж!D��s�!�_n�V����>y�e�⠹:TJ�����!,Ts����� �^�2�R.��ޑ�ih�v�fx�^�0y8'X�k(�ӊ��X�y?a�!���ྪ'�o'o��WS-f�`^��p�s���>�Vr�βVO�})yѧ� ]�5����*��~cB.i�E�����>��)�\y�8��s�*Zg�G"Ul�}�^пc��y����}�v�qy���a�F#b��
���nS�t� �m/>��/t��M�	�%[%�F*�y.�qV��-��,G���;�����3��A�֗�7߸ā�&
�;ڋzB��f�8<J8�������8��ax	3Sb�����]��g��IͿ����E���#�T� j���ZwLg֤�e�1~��vt���	y�����^?o�3��bI�1F��z�/-�2�Dwi�Z�r���SV0���h-iL�l����x�ͧM`��C�������%*�*@�� ��(�g��PG-/�)i'kdܶx��,p��m>!���訮lQ�;�p����qndwИ_[aqv�ABNn���uS�^�c��-O>�s��TUdx�du�y$X��/��R&��Zy���eѡ!�U��B���ʄ\kG)M�8��v���Y�5LqV�����/��;y�/�ct��>C�Ճ�OU(�C���	���}8֝O�O��B��
�;Ɓ�����k9��XS��4K#�7����=M�·�,�hm�2����¶sf����h��+�p�]���I"���)��O�1"��]����hݼ2�ҶΊ�K4���vi��J��c�!�_SrL���zlP�.�"���/#�w[�3(�����4��Z; �þ��2� ��d�,g42ut����qʅ�|����I�R�v�8��c-�O۝�i��ذՕ���$D��,���I��v�*�/�8S,�qx�٘~��aX�IvF>>�K��<�m���'�$�������L���9�n��$�F�A�n�]��Dқ�R�i�L�+���T{Gxh�a�b�1�	PPf�sR׋�^i�3��Wl�gkh�x2�������?��ѧ��4Ty}6T�ِ�q������ʞ)�M��]�����0��K����g�Hfk�x'V�ت?�)��y����>&���B�ñ!�����?��:�:��SM#`�*Obg-�홶/?7�8C�Y��b�X���yu��WR5��$��szO�@ߓ��Zl(��E�L
��e���Lv�6��[%:��.��MY��pwڌ�Q�K[�3奙ҵ%rw��l�DC(wo̕^����	�kփ�>��U�H�W�����P�8�pL����ӂH��6�_D����R�Vo�N�8
w�ZP��}�H�l���`hds��(t��9�����D���iڷ��V�̔�V�_u\��/K\�urB��핛�o�D?�O��XB1Q��6e�Ƿ��ďBA]��m��h꡼�Tj� D0-\�ލ��i�q�S�fI_]��ZyԎ��s�vz0��V��u5,C���HϽ�a6_�-"��\Y��\��YN��J�9��:hv�{T��c!�K��@)��;�j�V���!W�7�<�dX�G)k��"�� �J�<4}q�;�w��B0E��*e�·�׆�l�	2H7M5~��c_,밾钒�检"����K�_�F�@�>���9��*��z*���C!L��W�}\:�~Zu;���D� �흳���$��ng���)u� :2�{wVN�":��w�jNg�O�y�A:#ب�x�'+��1���A~6�!|9\m��'�?�]�lC,�B#��m���p�FWCk���I�j����D�K�9(^�L��w�,����@T!�9
M�_�T=fG�� S��x2��*YuՀCgt����o��?�HҮD9�y� ���ݍ�"�8��}�z�T��(�^*����;{�7��ZZ�Nl���4a�\ξ�`.��O�WcXUS�Mi�e؅Fj��\��B���_ ��9�e1��d��+�	��2��IWg����_>ѻyБ^#��/�[L���b���#.�1��>�[�����gT��b��o/6����&k�"dh���PrPR�c�x!�E��"X�C2�3��T9!=Ce���=�䏒_3l3f!�F��"�.i����\jD ����S�Ѩʄ7LI����UR�G	;���/<��j�!��?+�
� y�L�����I>�g1cԙ�+�t���n�Rk4�HEsL�Xp%�p�3�Ŭ� ��oi�-8��{v�9�Ъ��2L�ҁٕ���֘ʨX�� >@���l+�<�oo�]㲰V���F;��YѧWݚ�E]q���%��=�{�dW�>Б��9��AB���
�ᄯ�^N-Ҡo1{�1���h���G�X� �L��%=�J�+���+�ժ�z�E���	��� 7�~�ذ0sg0�F6 qb��9�L_�d7�dD�d���X�bkMJ`})L%��s�WFbe���.��M���l�Z}ή�w'����ND]��3m�,��O���%R��2�/)���V׆Z��`}��W�p-�ܧ���MU���g�����B�X�@��Cuw�į�bZ�xK������s=�s���O���q��g1�瓿4��, ez�H�Oh���@��wO��fCy"�/ꂨ{F"ѩuXX
�A����@!Ms	����&8O*h�Q`>��`�[�'�'[kϼO~qb+����,ј��V@ }�Xo���}�р�opV��~ؔR��N
���	�vy,������	I���B\B��*�xx�rX 5ԉ�JGO�r�m���Мp-,����L����;�����3�s��ekC̪-��w��#�]$ʄoT.���ҷA����(�X�-�*&z�O�0L�����Դ	۫�/�P�T�*8�%GhE�R��(�,�`	���҇4�=��4���&�����&�R��|:(<Kf��qA<E�We y�0[8Rz�������OX��@�Slߤ���'~�R����]��w7A�anQ���?���)�i�51_�A�zJ��(�M�y��k
��]RR俞�G�Cz깈��.+ܖ�:�Jwd�ۛ�D�e�?��@Z@<}L�~ßy(�k�GMd�j/W�a�w�Hh7��y��t�GI���[�ܦ��$Y�ݺV
	�;Yы�;���
��T.'�ι� �@L|�;��E
��3����[I��@��o�yv��5�EA8��J}\#���G��:!,���a���鑐�şv�k&IrNB��,���F��Ͳ���Iw8er�+��G����Zh<c���_U� ؏��D�s�����B�	�c�[�vKiNm��EX�����;$Ũj�!�������H�PQ�+��B�ᐻ}Y/���S���$3�ܚ]J����e4�4{���J*ό�7���	r�}#�$ej�U�G�-+B�>N��-��1�֣��LI	=��_�f��-&�e��wT	{������ɘ�� =O�P����:Z�裧�xAW�ne*3[��؜{�&�87N}��z$�㵓�4G��픶L�>�ǖ��[EY��t -���R��!�C�C��<*]ӯ�|�ٯ��߽�q����*, MR�m�y�e�r��-�/AW33�"󇄇��R���`�t0���ڂS��R{zH�L[W�Q��A"|6�]��DX�q�F�o���S��~���G{�sEp���8��,��W�	��Uʲ�?�J=���1�-�^"�����NWY���� �=��fl�HO�o��F1�H*x�7�1Fp�5⌻(wv�_Z���\��a��6���ro�fcAE���	���SbUl��g�Q�����'Cw\�ӳu$z��Uo���\�Z�M�x���*>�2p��������H
]7���88�͏}�~���L	�hP4����ê@Y��X@��Cx=m
�:ؙw^Mj�#����I4�L��.7�c����&}$��	�(�༝I"�16��)�a�|��%�a߂�0�7�Ȓ�i�����������"ረ2�bhn>
R鷋I�����};w*Zھvd�\ ���w�6@����ܦ���z�t&[��~z���`VL���8.��:��9�:x�����+H�*���o�,�-�Lj8�?T���Ɋ������wӢ�Iν���H�Teʫ�i��P��C�F�(������՝|��%�/����8j��#�S�M,��>�����z$=U�!E��ߞ=�9��"�E����#�<���^�TD l6���t�I����f '�W�|yو��K��w��Ԗ|��<�Z�w"o���p]�՗�(aj�ӋV�E�B��6ʵ���|�������V�_��_�ld�y�*��|\�SP�jѡq0s�km����ve�t����#�0�.ЋL�by����gx
<{<[HP����}�@G^��ũV?����ܶ4;K9�s�3RW��xF&-�:�3'��j�ӻT�k�HƦF�N����=�ߩ~���D�H�x��K��3�p8=ءXQ�2����=��®����uCao�"eD�p\S;�)��?�_��&�zϷ#���r�"eO=or.r��n>�Z��\Z$���w  �o����`��FV-Њ�l�l�����q��H)y�Z��<�C��8�е���C�7��7��D���͈��f?�d� �Ѹ!&�2�]��^�!�9�DZ���8��h���d�4~���!?��*���nr�{�9�.��h3f�x*�q�S���FƇv`k}Z�3-�x8z�������e�Q���s�c���b���߮ �B NT[\,3�@}5�g�'(�&'��듛�%�J��!_!���40퐵���%�|V��.��M4��^��ǿf���˭��#	�p��R^E�C��<�RJ�w�&�qG_P�*�I�XTu���ƙ!��w��H^��Kŏ�$B׏�~`�\q/�d6����`v �i~��*{�.+�|��C9[�|����ڣ�P�
nXT!T�]	F7�A�v�X����iǰ$w�mkR��ӥ����e#�`�6?�x��AM�l�}�/y"\g_� 
qޫl	��#��?����D��W"~�&F���N�k:J,�5 ��'���FO�g"OO"}WZ�"�_�&'R�8�>#A?%(���x22��`raw���{���`YT�����<�!��o&��ޥZl�j]��#��U>d3�J�x�W,s�p�a?3�h�%Em�(��B_����lqi
Ϣ&w`�l�o�[��9���T��7����IO�c�X��8.l��)k�2;���xoږ�:+.�b�a3OK�A<����*#cPv#q���::)�,Y%��k���$S�.`~D�>5�r��4#ծ^(��X�͋�bf��!�?�H��7J!�%�|͞�h��5Fg�_6x��!%¥��P]�NP������~���QJ/n�O��D��N���''���*گ��C	碔c��d�>��2_�|o}u��]�?0f�AL�?З��X�b��̿c[���3s�����a�m+����b��]�l�wgi]\�b��_�v��� y��g^̉tM�r�C���D(䚩_�&j�$W
˪���[E�ę��+"��Nl]@�݆BC:fJ���k�Gf�Ț�w��N�Wg'��5�b��	����uy�U@b��+X�7��a��	��	���6��-��s��b]�SI<鼭p�tqF�����L����$�۔����Yc��M���!���d�zmlP�!��d����#���"�$�O�������������<#�X�����ф��28R�Y֑n��ZKL���/��/a�,|'}���Щ�+��*����	R���������!���L��"VWզ�+f����9���t%#v3��a�	!:�E��YC�m!_q����Z�6�������۴fa��P��VQ�hT�*
��K��u�5��v��)uw�M����*C�4�$B��ZVi������$��)����q�q�	��l�A�Q1�n�i+�KI[�{�3#W�;�Q��w�X�խZ�C![�<#�O����3�q[.U�R��K��OP�¤�h���m�F����tU��~�B�,)xH�Pd��a"$ q;*��(W΂r�Q{	��5%�K���o�n^S�q���4�-?>#�~��Lª�بw��2ꔔ��PCS{��X��VG�T�jO0���L�ĞN܅4�K��Q*'1�h"-6��`eJ��a��ih����������z�y~��3Di�U2Z�.��Akؽ2�GAχ��K_q�~�"2�=>��}:�9K���d-V�zj�Y��FR�����SUڀ��4Ռ��M���$�Amg.?��������ūT����?��5�%��Pd��}����Ϫ%����B��5�N r�����6%��u��6���wf>��nV�:���L��HV���ڜʌ��!q�(�E�q� ���i��bl�_�Sc����o�v�C". �h|ý (2�(��+.3K'�s�������.�6ӿ����|���k�"��,�p%b󿨆���k��黼ׁR^b0��ˡ4�vP%���A'��?�1��34F`\ZZ|o7t�	*�?��Lqٰ�Ѽ:w�m9Ss�cx4�∺L��Asî?D��'+��.�9��-�K�E�6�i2����:�e��tV�=�ԍ�[H}G3}"/ns0 �?��>�ly]�j��0V��E�6I�h;�_���S��QX	�vs�eH�H���1®ru}ϩ�y�!z���iC����֥�g'&�! ��*��fGb��6h�[m��[�VnD���/=޿4
����%��3�v��eW�q(�����f��2��j&���I�n]�r�a��M9��\�*z�$]R?	M��vv�ф��u�>?}��251���1�`�GG�:O�=SQ:wdȤ�S�\��yw�jm�_d�����&i.�	�6�O�P�3n`˿_O��� ��@�9�L�F=�M���:�6�B��f�1y�4����V"��l��²WU�=��2�կ��/aMҲ|���;7��QC����z
�Ң�N��b�*�]܎�m��".�r.�MU�訫��QzK�"i�ͅ0���	S��E�ȃ���/������� I�.C�<b2] $�Zƻ4����� ��obm��dcseA�X��4����&S������y}�^{�F�o+��I!��@�r��{FJ7����`��y��xDL	���Kդƾ��\ʢ[�3����k��c�;���6HzX[]]y EUe4y�8�uq�h�������W�-��K��=�閸9D���q��0�"W∕���,_dJP�1��"������LA[�h�xA�-ڛau���>7�ո��%�?aD323�2��`;�]���nҸ�#9�.%�pGiYl�j�qn�&lć&q~Yh0��S���.����=Q��8��է	�a��v%8g�U��w(쨴ȥڏ��4����Bͪ:OkC���x�"�a1$C�ņ������Y�	p�^7"q����ۋ�������( ��/q�qTڷ���0�